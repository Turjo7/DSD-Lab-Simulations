CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 476 52 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 P5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43544.5 0
0
13 Logic Switch~
5 417 50 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 P4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43544.5 0
0
13 Logic Switch~
5 89 97 0 1 11
0 2
0
0 0 21360 0
2 0V
-7 -12 7 -4
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
43544.5 0
0
13 Logic Switch~
5 191 103 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -17 8 -9
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
43544.5 0
0
13 Logic Switch~
5 341 49 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 P3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43544.5 0
0
13 Logic Switch~
5 271 49 0 1 11
0 8
0
0 0 21360 0
2 0V
-4 -16 10 -8
2 P2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
43544.5 0
0
13 Logic Switch~
5 198 51 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 P1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8901 0 0
2
43544.5 0
0
13 Logic Switch~
5 486 296 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7361 0 0
2
43544.5 0
0
13 Logic Switch~
5 261 219 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4747 0 0
2
43544.5 0
0
8 2-In OR~
219 359 371 0 3 22
0 4 3 18
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
972 0 0
2
43544.5 0
0
9 Inverter~
13 71 361 0 2 22
0 2 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3472 0 0
2
43544.5 0
0
8 3-In OR~
219 304 158 0 4 22
0 9 12 7 10
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 3 0
1 U
9998 0 0
2
43544.5 0
0
9 2-In AND~
219 177 369 0 3 22
0 6 5 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3536 0 0
2
43544.5 0
0
9 2-In AND~
219 178 307 0 3 22
0 2 11 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
4597 0 0
2
43544.5 0
0
9 2-In AND~
219 173 242 0 3 22
0 14 13 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3835 0 0
2
43544.5 0
0
6 74136~
219 123 193 0 3 22
0 2 15 14
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3670 0 0
2
43544.5 0
0
8 3-In OR~
219 296 334 0 4 22
0 9 8 7 4
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
5616 0 0
2
43544.5 0
0
14 Logic Display~
6 648 159 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9323 0 0
2
43544.5 0
0
7 Pulser~
4 321 228 0 11 12
0 19 21 20 22 0 0 5 5 -1
7 1
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
317 0 0
2
43544.5 0
0
6 JK RN~
219 516 226 0 6 22
0 10 20 18 16 23 17
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
3108 0 0
2
43544.5 0
0
24
1 1 2 0 0 4096 0 3 16 0 0 3
101 97
101 184
107 184
3 2 3 0 0 4224 0 13 10 0 0 4
198 369
329 369
329 380
346 380
4 1 4 0 0 4224 0 17 10 0 0 3
329 334
329 362
346 362
1 2 5 0 0 12416 0 1 13 0 0 6
488 52
721 52
721 423
135 423
135 378
153 378
2 1 6 0 0 8320 0 11 13 0 0 3
92 361
92 360
153 360
0 1 2 0 0 0 0 0 11 13 0 4
91 298
30 298
30 361
56 361
0 3 7 0 0 8192 0 0 17 11 0 3
221 307
221 343
283 343
1 2 8 0 0 12416 0 6 17 0 0 5
283 49
283 94
229 94
229 334
284 334
0 1 9 0 0 8320 0 0 17 15 0 4
212 242
259 242
259 325
283 325
4 0 10 0 0 4096 0 12 0 0 22 4
337 158
371 158
371 181
401 181
3 3 7 0 0 8320 0 14 12 0 0 5
199 307
221 307
221 178
291 178
291 167
1 2 11 0 0 8320 0 2 14 0 0 5
429 50
429 15
53 15
53 316
154 316
0 1 2 0 0 8320 0 0 14 1 0 4
101 183
91 183
91 298
154 298
1 2 12 0 0 8320 0 5 12 0 0 5
353 49
353 103
263 103
263 158
292 158
3 1 9 0 0 0 0 15 12 0 0 6
194 242
212 242
212 168
283 168
283 149
291 149
1 2 13 0 0 12416 0 7 15 0 0 5
210 51
210 71
41 71
41 251
149 251
3 1 14 0 0 8320 0 16 15 0 0 5
156 193
156 215
133 215
133 233
149 233
1 2 15 0 0 8320 0 4 16 0 0 5
203 103
203 126
81 126
81 202
107 202
1 4 16 0 0 8320 0 8 20 0 0 3
498 296
516 296
516 257
6 1 17 0 0 4224 0 20 18 0 0 3
540 209
648 209
648 177
3 3 18 0 0 8320 0 10 20 0 0 6
392 371
397 371
397 250
455 250
455 227
492 227
0 1 10 0 0 4224 0 0 20 0 0 4
398 181
455 181
455 209
492 209
1 1 19 0 0 4224 0 9 19 0 0 2
273 219
297 219
3 2 20 0 0 12416 0 19 20 0 0 4
345 219
357 219
357 218
485 218
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
