CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
220 10 30 110 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 921 179 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3536 0 0
2
43495.5 0
0
13 Logic Switch~
5 388 66 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4597 0 0
2
43495.5 0
0
13 Logic Switch~
5 473 65 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3835 0 0
2
43495.5 0
0
13 Logic Switch~
5 977 187 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3670 0 0
2
43495.5 0
0
13 Logic Switch~
5 1042 186 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5616 0 0
2
43495.5 0
0
7 Ground~
168 531 323 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9323 0 0
2
43495.5 0
0
2 +V
167 233 234 0 1 3
0 7
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
317 0 0
2
43495.5 0
0
5 4049~
219 307 139 0 2 22
0 3 5
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
3108 0 0
2
43495.5 0
0
5 4049~
219 643 36 0 2 22
0 4 6
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
4299 0 0
2
43495.5 0
0
14 Logic Display~
6 1143 98 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9672 0 0
2
43495.5 0
0
14 Logic Display~
6 1200 103 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7876 0 0
2
43495.5 0
0
7 Ground~
168 812 292 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6369 0 0
2
43495.5 0
0
7 74LS151
20 642 406 0 14 29
0 7 2 4 4 4 2 5 3 2
10 11 12 8 13
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
9172 0 0
2
43495.5 0
0
7 74LS151
20 642 185 0 14 29
0 7 2 3 3 2 3 6 4 2
10 11 12 9 14
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
7100 0 0
2
43495.5 0
0
28
0 3 3 0 0 8192 0 0 14 10 0 3
347 82
347 176
610 176
0 3 4 0 0 4096 0 0 13 18 0 3
546 65
546 397
610 397
0 4 4 0 0 4096 0 0 13 18 0 3
509 65
509 406
610 406
0 4 3 0 0 0 0 0 14 17 0 4
421 109
541 109
541 185
610 185
0 5 2 0 0 8192 0 0 14 14 0 4
531 295
588 295
588 194
610 194
0 5 4 0 0 4224 0 0 13 18 0 3
493 65
493 415
610 415
0 6 2 0 0 8192 0 0 13 14 0 4
531 307
563 307
563 424
610 424
0 6 3 0 0 0 0 0 14 17 0 4
421 213
550 213
550 203
610 203
2 7 5 0 0 8320 0 8 13 0 0 4
328 139
472 139
472 433
610 433
0 1 3 0 0 0 0 0 8 17 0 4
421 82
275 82
275 139
292 139
2 7 6 0 0 12416 0 9 14 0 0 6
664 36
691 36
691 123
585 123
585 212
610 212
0 1 4 0 0 0 0 0 9 18 0 3
524 65
524 36
628 36
0 2 2 0 0 0 0 0 13 14 0 4
531 283
600 283
600 388
610 388
1 2 2 0 0 4224 0 6 14 0 0 3
531 317
531 167
610 167
0 1 7 0 0 8320 0 0 13 16 0 3
272 252
272 379
610 379
1 1 7 0 0 0 0 7 14 0 0 5
233 243
233 252
522 252
522 158
610 158
1 8 3 0 0 8320 0 2 13 0 0 4
400 66
421 66
421 442
610 442
1 8 4 0 0 128 0 3 14 0 0 4
485 65
558 65
558 221
610 221
13 1 8 0 0 4224 0 13 10 0 0 3
674 433
1143 433
1143 116
13 1 9 0 0 4224 0 14 11 0 0 3
674 212
1200 212
1200 121
0 9 2 0 0 0 0 0 13 22 0 4
812 271
709 271
709 379
680 379
1 9 2 0 0 128 0 12 14 0 0 3
812 286
812 158
680 158
0 10 10 0 0 8320 0 0 13 26 0 3
1027 256
1027 388
674 388
0 11 11 0 0 8192 0 0 13 27 0 3
953 237
953 397
674 397
0 12 12 0 0 4096 0 0 13 28 0 3
873 199
873 406
674 406
1 10 10 0 0 0 0 5 14 0 0 6
1054 186
1078 186
1078 256
786 256
786 167
674 167
1 11 11 0 0 12416 0 4 14 0 0 6
989 187
1001 187
1001 237
716 237
716 176
674 176
1 12 12 0 0 20608 0 1 14 0 0 8
933 179
944 179
944 186
920 186
920 199
696 199
696 185
674 185
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
