CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 80 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 100 28 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7346 0 0
2
43490.9 0
0
13 Logic Switch~
5 26 29 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8577 0 0
2
43490.9 0
0
13 Logic Switch~
5 137 1429 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3372 0 0
2
43490.9 0
0
13 Logic Switch~
5 96 1431 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3741 0 0
2
43490.9 0
0
13 Logic Switch~
5 61 1432 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5813 0 0
2
43490.9 0
0
2 +V
167 1035 408 0 1 3
0 3
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3213 0 0
2
43490.9 0
0
7 Ground~
168 1009 333 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3694 0 0
2
43490.9 0
0
5 4049~
219 70 91 0 2 22
0 5 6
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U12E
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 12 0
1 U
4327 0 0
2
43490.9 0
0
5 4049~
219 22 96 0 2 22
0 4 7
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U12D
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 12 0
1 U
8800 0 0
2
43490.9 0
0
5 4049~
219 161 1324 0 2 22
0 8 11
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U12C
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 12 0
1 U
3406 0 0
2
43490.9 0
0
5 4049~
219 99 1324 0 2 22
0 9 12
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U12B
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 12 0
1 U
6455 0 0
2
43490.9 0
0
5 4049~
219 45 1325 0 2 22
0 10 14
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U12A
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 12 0
1 U
9319 0 0
2
43490.9 0
0
14 Logic Display~
6 872 55 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3172 0 0
2
43490.9 0
0
14 Logic Display~
6 810 58 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
38 0 0
2
43490.9 0
0
5 4071~
219 642 927 0 3 22
0 18 17 15
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 11 0
1 U
376 0 0
2
43490.9 0
0
5 4071~
219 633 221 0 3 22
0 28 27 16
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 11 0
1 U
6666 0 0
2
43490.9 0
0
8 4-In OR~
219 485 1045 0 5 22
0 22 21 20 19 17
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U10B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
9365 0 0
2
43490.9 0
0
8 4-In OR~
219 487 824 0 5 22
0 26 25 24 23 18
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U10A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
3251 0 0
2
43490.9 0
0
8 4-In OR~
219 481 359 0 5 22
0 32 31 30 29 27
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U9B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 9 0
1 U
5481 0 0
2
43490.9 0
0
8 4-In OR~
219 471 114 0 5 22
0 36 35 34 33 28
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U9A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 9 0
1 U
7788 0 0
2
43490.9 0
0
5 4082~
219 286 1179 0 5 22
0 3 10 9 8 19
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 8 0
1 U
3273 0 0
2
43490.9 0
0
5 4082~
219 287 1115 0 5 22
0 2 10 9 11 20
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 8 0
1 U
3761 0 0
2
43490.9 0
0
5 4082~
219 289 1049 0 5 22
0 4 10 12 8 21
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U7B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 7 0
1 U
3226 0 0
2
43490.9 0
0
5 4082~
219 290 985 0 5 22
0 4 10 12 11 22
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U7A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
4244 0 0
2
43490.9 0
0
5 4082~
219 290 916 0 5 22
0 2 14 9 8 23
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U6B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 6 0
1 U
5225 0 0
2
43490.9 0
0
5 4082~
219 292 845 0 5 22
0 4 14 9 11 24
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U6A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
768 0 0
2
43490.9 0
0
5 4082~
219 291 774 0 5 22
0 6 14 12 8 25
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
5735 0 0
2
43490.9 0
0
5 4082~
219 292 692 0 5 22
0 5 14 12 11 26
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
5881 0 0
2
43490.9 0
0
5 4082~
219 297 528 0 5 22
0 3 10 9 8 29
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
3275 0 0
2
43490.9 0
0
5 4082~
219 299 456 0 5 22
0 2 10 9 11 30
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
4203 0 0
2
43490.9 0
0
5 4082~
219 302 386 0 5 22
0 5 13 12 8 31
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
3440 0 0
2
43490.9 0
0
5 4082~
219 303 320 0 5 22
0 5 10 12 11 32
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
9102 0 0
2
43490.9 0
0
5 4082~
219 308 60 0 5 22
0 4 14 12 11 36
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
5586 0 0
2
43490.9 0
0
5 4082~
219 305 253 0 5 22
0 5 14 9 8 33
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
525 0 0
2
43490.9 0
0
5 4082~
219 305 193 0 5 22
0 2 14 9 11 34
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
6206 0 0
2
43490.9 0
0
5 4082~
219 306 129 0 5 22
0 7 14 12 8 35
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 1 0
1 U
3418 0 0
2
43490.9 0
0
91
0 1 3 0 0 8320 0 0 21 2 0 5
1010 497
1010 1144
221 1144
221 1166
262 1166
1 1 3 0 0 0 0 6 29 0 0 5
1035 417
1035 497
253 497
253 515
273 515
0 1 2 0 0 4224 0 0 22 4 0 5
960 314
960 1078
250 1078
250 1102
263 1102
0 1 2 0 0 0 0 0 30 11 0 6
1009 314
642 314
642 419
265 419
265 443
275 443
0 1 4 0 0 4224 0 0 23 18 0 3
235 47
235 1036
265 1036
0 1 5 0 0 8192 0 0 31 17 0 3
132 371
132 373
278 373
0 1 5 0 0 8192 0 0 32 10 0 4
123 19
189 19
189 307
279 307
0 1 4 0 0 128 0 0 24 18 0 7
44 29
44 12
682 12
682 951
236 951
236 972
266 972
0 1 2 0 0 0 0 0 25 11 0 6
1009 285
711 285
711 872
250 872
250 903
266 903
0 1 5 0 0 0 0 0 34 17 0 5
123 28
123 5
200 5
200 240
281 240
1 1 2 0 0 128 0 7 35 0 0 7
1009 327
1009 259
404 259
404 159
272 159
272 180
281 180
0 1 4 0 0 128 0 0 26 16 0 6
25 63
7 63
7 814
262 814
262 832
268 832
2 1 6 0 0 4224 0 8 27 0 0 3
73 109
73 761
267 761
0 1 5 0 0 0 0 0 8 17 0 3
132 38
73 38
73 73
2 1 7 0 0 4224 0 9 36 0 0 4
25 114
273 114
273 116
282 116
0 1 4 0 0 0 0 0 9 18 0 3
67 37
25 37
25 78
1 1 5 0 0 8320 0 1 28 0 0 6
112 28
132 28
132 626
259 626
259 679
268 679
1 1 4 0 0 128 0 2 33 0 0 4
38 29
67 29
67 47
284 47
0 4 8 0 0 4096 0 0 21 56 0 4
151 1198
258 1198
258 1193
262 1193
0 4 8 0 0 8192 0 0 29 56 0 3
151 543
151 542
273 542
0 3 9 0 0 8192 0 0 21 52 0 3
83 1185
83 1184
262 1184
0 3 9 0 0 8192 0 0 29 52 0 3
83 532
83 533
273 533
0 2 10 0 0 4096 0 0 21 42 0 4
17 1178
225 1178
225 1175
262 1175
0 2 10 0 0 8192 0 0 29 42 0 3
17 523
17 524
273 524
0 4 11 0 0 8192 0 0 22 64 0 3
164 1130
164 1129
263 1129
0 4 11 0 0 4096 0 0 30 64 0 4
164 474
271 474
271 470
275 470
0 3 9 0 0 0 0 0 22 52 0 3
83 1121
83 1120
263 1120
0 3 9 0 0 8192 0 0 30 52 0 3
83 463
83 461
275 461
0 2 10 0 0 0 0 0 22 42 0 3
17 1110
17 1111
263 1111
0 2 10 0 0 8192 0 0 30 42 0 3
17 451
17 452
275 452
0 4 8 0 0 0 0 0 23 56 0 3
151 1061
151 1063
265 1063
0 4 8 0 0 0 0 0 31 56 0 4
151 405
271 405
271 400
278 400
0 3 12 0 0 8192 0 0 23 65 0 3
102 1055
102 1054
265 1054
0 3 12 0 0 0 0 0 31 65 0 4
102 394
232 394
232 391
278 391
0 2 10 0 0 0 0 0 23 42 0 3
17 1043
17 1045
265 1045
0 2 13 0 0 4224 0 0 31 0 0 2
20 382
278 382
0 4 11 0 0 0 0 0 24 64 0 3
164 1000
164 999
266 999
0 4 11 0 0 4096 0 0 32 64 0 4
164 338
273 338
273 334
279 334
0 3 12 0 0 8192 0 0 24 65 0 3
102 989
102 990
266 990
0 3 12 0 0 8192 0 0 32 65 0 3
102 326
102 325
279 325
0 2 10 0 0 0 0 0 24 42 0 3
17 982
17 981
266 981
0 2 10 0 0 8320 0 0 32 69 0 4
73 1361
17 1361
17 316
279 316
0 4 8 0 0 0 0 0 25 56 0 2
151 930
266 930
0 4 8 0 0 8192 0 0 34 56 0 3
151 268
151 267
281 267
0 3 9 0 0 0 0 0 25 52 0 3
83 922
83 921
266 921
0 3 9 0 0 8192 0 0 34 52 0 3
83 257
83 258
281 258
0 2 14 0 0 8192 0 0 25 66 0 3
48 911
48 912
266 912
0 2 14 0 0 4096 0 0 34 66 0 2
48 249
281 249
0 4 11 0 0 0 0 0 26 64 0 3
164 860
164 859
268 859
0 4 11 0 0 8192 0 0 35 64 0 3
164 206
164 207
281 207
0 3 9 0 0 0 0 0 26 52 0 2
83 850
268 850
0 3 9 0 0 8320 0 0 35 68 0 4
102 1345
83 1345
83 198
281 198
0 2 14 0 0 0 0 0 26 66 0 4
48 832
244 832
244 841
268 841
0 2 14 0 0 0 0 0 35 66 0 4
48 193
254 193
254 189
281 189
0 4 8 0 0 0 0 0 27 56 0 3
151 787
151 788
267 788
0 4 8 0 0 8320 0 0 36 67 0 6
164 1365
151 1365
151 151
277 151
277 143
282 143
0 3 12 0 0 0 0 0 27 65 0 3
102 781
102 779
267 779
0 2 14 0 0 0 0 0 27 66 0 3
48 769
48 770
267 770
0 3 12 0 0 0 0 0 36 65 0 4
102 141
234 141
234 134
282 134
0 2 14 0 0 8192 0 0 36 66 0 3
48 124
48 125
282 125
0 4 11 0 0 0 0 0 28 64 0 2
164 706
268 706
0 3 12 0 0 0 0 0 28 65 0 3
102 694
102 697
268 697
0 2 14 0 0 0 0 0 28 66 0 4
48 672
223 672
223 688
268 688
2 4 11 0 0 4224 0 10 33 0 0 3
164 1306
164 74
284 74
2 3 12 0 0 4224 0 11 33 0 0 3
102 1306
102 65
284 65
2 2 14 0 0 4224 0 12 33 0 0 3
48 1307
48 56
284 56
1 1 8 0 0 0 0 3 10 0 0 3
149 1429
164 1429
164 1342
1 1 9 0 0 0 0 4 11 0 0 5
108 1431
119 1431
119 1350
102 1350
102 1342
1 1 10 0 0 0 0 5 12 0 0 4
73 1432
73 1349
48 1349
48 1343
3 1 15 0 0 8320 0 15 13 0 0 5
675 927
867 927
867 82
872 82
872 73
3 1 16 0 0 8320 0 16 14 0 0 3
666 221
810 221
810 76
5 2 17 0 0 8320 0 17 15 0 0 4
518 1045
600 1045
600 936
629 936
5 1 18 0 0 8320 0 18 15 0 0 4
520 824
599 824
599 918
629 918
5 4 19 0 0 4224 0 21 17 0 0 4
307 1179
453 1179
453 1059
468 1059
5 3 20 0 0 4224 0 22 17 0 0 4
308 1115
439 1115
439 1050
468 1050
5 2 21 0 0 4224 0 23 17 0 0 4
310 1049
418 1049
418 1041
468 1041
5 1 22 0 0 4224 0 24 17 0 0 4
311 985
452 985
452 1032
468 1032
5 4 23 0 0 4224 0 25 18 0 0 6
311 916
418 916
418 859
447 859
447 838
470 838
5 3 24 0 0 4224 0 26 18 0 0 4
313 845
417 845
417 829
470 829
5 2 25 0 0 4224 0 27 18 0 0 4
312 774
446 774
446 820
470 820
5 1 26 0 0 4224 0 28 18 0 0 4
313 692
460 692
460 811
470 811
5 2 27 0 0 8320 0 19 16 0 0 4
514 359
603 359
603 230
620 230
5 1 28 0 0 4224 0 20 16 0 0 4
504 114
602 114
602 212
620 212
5 4 29 0 0 8320 0 29 19 0 0 4
318 528
356 528
356 373
464 373
5 3 30 0 0 12416 0 30 19 0 0 4
320 456
347 456
347 364
464 364
5 2 31 0 0 12416 0 31 19 0 0 4
323 386
336 386
336 355
464 355
5 1 32 0 0 4224 0 32 19 0 0 4
324 320
444 320
444 346
464 346
5 4 33 0 0 8320 0 34 20 0 0 4
326 253
356 253
356 128
454 128
5 3 34 0 0 12416 0 35 20 0 0 4
326 193
346 193
346 119
454 119
5 2 35 0 0 12416 0 36 20 0 0 6
327 129
336 129
336 77
432 77
432 110
454 110
5 1 36 0 0 4224 0 33 20 0 0 4
329 60
443 60
443 101
454 101
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
856 4 893 28
866 12 882 28
2 F1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
788 8 825 32
798 16 814 32
2 F0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
