CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 40 380 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 41 288 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 38 179 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 38 75 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 256 575 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 187 575 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89878e-315 0
0
5 4049~
219 272 490 0 2 22
0 2 4
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U4B
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 4 0
1 U
8901 0 0
2
5.89878e-315 0
0
5 4049~
219 190 490 0 2 22
0 3 5
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U4A
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
7361 0 0
2
5.89878e-315 0
0
14 Logic Display~
6 1024 229 0 1 2
10 10
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.89878e-315 0
0
8 4-In OR~
219 805 230 0 5 22
0 14 13 12 11 10
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
972 0 0
2
5.89878e-315 0
0
5 7415~
219 416 412 0 4 22
0 6 3 2 11
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 2 0
1 U
3472 0 0
2
5.89878e-315 0
0
5 7415~
219 418 303 0 4 22
0 7 3 4 12
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 1 0
1 U
9998 0 0
2
5.89878e-315 0
0
5 7415~
219 419 191 0 4 22
0 8 5 2 13
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
3536 0 0
2
5.89878e-315 0
0
5 7415~
219 420 98 0 4 22
0 9 5 4 14
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
4597 0 0
2
5.89878e-315 0
0
19
0 3 2 0 0 4096 0 0 11 5 0 4
241 426
381 426
381 421
392 421
0 2 3 0 0 4096 0 0 11 4 0 4
144 407
381 407
381 412
392 412
0 3 4 0 0 4096 0 0 12 7 0 3
275 315
394 315
394 312
0 2 3 0 0 12416 0 0 12 10 0 4
199 533
144 533
144 303
394 303
0 3 2 0 0 8320 0 0 13 9 0 4
311 530
241 530
241 200
395 200
0 2 5 0 0 4096 0 0 13 8 0 2
193 191
395 191
2 3 4 0 0 4224 0 7 14 0 0 3
275 472
275 107
396 107
2 2 5 0 0 4224 0 8 14 0 0 3
193 472
193 98
396 98
1 1 2 0 0 0 0 5 7 0 0 5
268 575
311 575
311 516
275 516
275 508
1 1 3 0 0 0 0 6 8 0 0 4
199 575
199 515
193 515
193 508
1 1 6 0 0 4224 0 1 11 0 0 4
52 380
382 380
382 403
392 403
1 1 7 0 0 4224 0 2 12 0 0 4
53 288
383 288
383 294
394 294
1 1 8 0 0 8320 0 3 13 0 0 3
50 179
50 182
395 182
1 1 9 0 0 4224 0 4 14 0 0 4
50 75
384 75
384 89
396 89
5 1 10 0 0 8320 0 10 9 0 0 3
838 230
838 233
1008 233
4 4 11 0 0 4224 0 11 10 0 0 4
437 412
769 412
769 244
788 244
4 3 12 0 0 4224 0 12 10 0 0 4
439 303
755 303
755 235
788 235
4 2 13 0 0 4224 0 13 10 0 0 4
440 191
755 191
755 226
788 226
4 1 14 0 0 4224 0 14 10 0 0 4
441 98
769 98
769 217
788 217
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
