CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
60 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
81
13 Logic Switch~
5 721 247 0 1 11
0 68
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6891 0 0
2
43514 0
0
13 Logic Switch~
5 446 253 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5407 0 0
2
43514 0
0
13 Logic Switch~
5 546 255 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7349 0 0
2
43514 0
0
13 Logic Switch~
5 626 253 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3919 0 0
2
43514 0
0
13 Logic Switch~
5 231 111 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9747 0 0
2
43514 0
0
13 Logic Switch~
5 313 112 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5310 0 0
2
43514 0
0
13 Logic Switch~
5 386 113 0 10 11
0 52 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4318 0 0
2
43514 0
0
13 Logic Switch~
5 478 109 0 10 11
0 72 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3917 0 0
2
43514 0
0
13 Logic Switch~
5 228 45 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7930 0 0
2
43514 0
0
13 Logic Switch~
5 316 46 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6128 0 0
2
43514 0
0
13 Logic Switch~
5 399 45 0 10 11
0 56 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7346 0 0
2
43514 0
0
13 Logic Switch~
5 476 42 0 10 11
0 74 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8577 0 0
2
43514 0
0
14 Logic Display~
6 717 62 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3372 0 0
2
43514 0
0
5 4071~
219 2358 2971 0 3 22
0 4 3 2
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U13D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 13 0
1 U
3741 0 0
2
43514 0
0
5 4081~
219 2271 3010 0 3 22
0 5 6 3
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U16D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 16 0
1 U
5813 0 0
2
43514 0
0
5 4081~
219 2299 2909 0 3 22
0 8 7 4
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U16C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 16 0
1 U
3213 0 0
2
43514 0
0
5 4030~
219 2220 2842 0 3 22
0 5 6 8
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U14D
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 14 0
1 U
3694 0 0
2
43514 0
0
5 4030~
219 2086 3161 0 3 22
0 10 7 9
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U14C
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 14 0
1 U
4327 0 0
2
43514 0
0
5 4030~
219 2028 3061 0 3 22
0 5 6 10
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U14B
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 14 0
1 U
8800 0 0
2
43514 0
0
5 4049~
219 1429 3164 0 2 22
0 11 12
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11F
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 11 0
1 U
3406 0 0
2
43514 0
0
5 4081~
219 1645 3181 0 3 22
0 12 13 7
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U16B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 16 0
1 U
6455 0 0
2
43514 0
0
5 4049~
219 1405 2936 0 2 22
0 16 17
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11E
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 11 0
1 U
9319 0 0
2
43514 0
0
5 4071~
219 1597 2981 0 3 22
0 19 18 6
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U13C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 13 0
1 U
3172 0 0
2
43514 0
0
5 4081~
219 1509 3021 0 3 22
0 14 16 18
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U16A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 16 0
1 U
38 0 0
2
43514 0
0
5 4081~
219 1507 2953 0 3 22
0 17 15 19
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U12D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 12 0
1 U
376 0 0
2
43514 0
0
5 4071~
219 1411 2600 0 3 22
0 21 20 5
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U13B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 13 0
1 U
6666 0 0
2
43514 0
0
5 4049~
219 1037 2591 0 2 22
0 14 22
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11D
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 11 0
1 U
9365 0 0
2
43514 0
0
5 4073~
219 1255 2572 0 4 22
0 23 11 22 21
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U15A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 15 0
1 U
3251 0 0
2
43514 0
0
5 4030~
219 1159 2536 0 3 22
0 16 15 23
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U14A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 14 0
1 U
5481 0 0
2
43514 0
0
5 4071~
219 1432 2368 0 3 22
0 25 24 13
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U13A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 13 0
1 U
7788 0 0
2
43514 0
0
5 4081~
219 1361 2409 0 3 22
0 27 26 24
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U12C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 12 0
1 U
3273 0 0
2
43514 0
0
5 4081~
219 1357 2344 0 3 22
0 29 28 25
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U12B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 12 0
1 U
3761 0 0
2
43514 0
0
5 4030~
219 1237 2332 0 3 22
0 27 26 29
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U10D
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 10 0
1 U
3226 0 0
2
43514 0
0
5 4030~
219 1212 2072 0 3 22
0 31 28 30
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U10C
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 10 0
1 U
4244 0 0
2
43514 0
0
5 4030~
219 1166 1973 0 3 22
0 27 26 31
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U10B
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 10 0
1 U
5225 0 0
2
43514 0
0
5 4049~
219 727 2266 0 2 22
0 11 32
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11C
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 11 0
1 U
768 0 0
2
43514 0
0
5 4081~
219 906 2261 0 3 22
0 33 32 28
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U12A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 12 0
1 U
5735 0 0
2
43514 0
0
5 4049~
219 664 2069 0 2 22
0 34 35
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11B
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 11 0
1 U
5881 0 0
2
43514 0
0
5 4071~
219 909 2105 0 3 22
0 37 36 26
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U8D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 8 0
1 U
3275 0 0
2
43514 0
0
5 4081~
219 778 2150 0 3 22
0 14 34 36
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 9 0
1 U
4203 0 0
2
43514 0
0
5 4081~
219 776 2057 0 3 22
0 15 35 37
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 9 0
1 U
3440 0 0
2
43514 0
0
5 4071~
219 967 1899 0 3 22
0 39 38 27
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 8 0
1 U
9102 0 0
2
43514 0
0
5 4049~
219 594 1925 0 2 22
0 14 40
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 11 0
1 U
5586 0 0
2
43514 0
0
5 4073~
219 833 1847 0 4 22
0 41 11 40 39
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 2 0
1 U
525 0 0
2
43514 0
0
5 4030~
219 723 1825 0 3 22
0 15 34 41
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U10A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 10 0
1 U
6206 0 0
2
43514 0
0
5 4071~
219 1532 1554 0 3 22
0 43 42 33
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 8 0
1 U
3418 0 0
2
43514 0
0
5 4081~
219 1450 1615 0 3 22
0 45 44 42
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 9 0
1 U
9312 0 0
2
43514 0
0
5 4081~
219 1452 1511 0 3 22
0 47 46 43
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 9 0
1 U
7419 0 0
2
43514 0
0
5 4030~
219 1357 1483 0 3 22
0 45 44 47
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U7D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 7 0
1 U
472 0 0
2
43514 0
0
5 4030~
219 1243 1421 0 3 22
0 49 46 48
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U7C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 7 0
1 U
4714 0 0
2
43514 0
0
5 4030~
219 1201 1340 0 3 22
0 45 44 49
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U7B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
9386 0 0
2
43514 0
0
5 4049~
219 653 1642 0 2 22
0 11 50
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
7610 0 0
2
43514 0
0
5 4081~
219 893 1626 0 3 22
0 51 50 46
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 6 0
1 U
3482 0 0
2
43514 0
0
5 4049~
219 688 1411 0 2 22
0 52 53
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
3608 0 0
2
43514 0
0
5 4071~
219 984 1460 0 3 22
0 55 54 44
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 8 0
1 U
6397 0 0
2
43514 0
0
5 4081~
219 904 1504 0 3 22
0 14 52 54
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 6 0
1 U
3967 0 0
2
43514 0
0
5 4081~
219 902 1423 0 3 22
0 53 15 55
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
8621 0 0
2
43514 0
0
5 4071~
219 1072 1269 0 3 22
0 57 56 45
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
8901 0 0
2
43514 0
0
5 4049~
219 742 1279 0 2 22
0 14 58
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
7385 0 0
2
43514 0
0
5 4073~
219 988 1258 0 4 22
0 59 11 58 57
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
6519 0 0
2
43514 0
0
5 4030~
219 843 1227 0 3 22
0 52 15 59
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U7A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
552 0 0
2
43514 0
0
5 4071~
219 1404 886 0 3 22
0 61 60 51
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
5551 0 0
2
43514 0
0
5 4081~
219 1324 930 0 3 22
0 63 62 60
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
8715 0 0
2
43514 0
0
5 4081~
219 1314 847 0 3 22
0 65 64 61
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
9763 0 0
2
43514 0
0
5 4030~
219 1180 814 0 3 22
0 63 62 65
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
8443 0 0
2
43514 0
0
5 4030~
219 1193 1045 0 3 22
0 67 64 66
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
3719 0 0
2
43514 0
0
5 4030~
219 1135 974 0 3 22
0 63 62 67
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
8671 0 0
2
43514 0
0
5 4049~
219 781 1027 0 2 22
0 11 69
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
7168 0 0
2
43514 0
0
5 4081~
219 948 1036 0 3 22
0 69 68 64
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
49 0 0
2
43514 0
0
5 4049~
219 766 903 0 2 22
0 72 73
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
6536 0 0
2
43514 0
0
5 4071~
219 1053 872 0 3 22
0 71 70 62
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
3931 0 0
2
43514 0
0
5 4081~
219 944 915 0 3 22
0 73 15 70
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
4390 0 0
2
43514 0
0
5 4081~
219 940 835 0 3 22
0 72 14 71
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
3242 0 0
2
43514 0
0
5 4071~
219 1046 726 0 3 22
0 75 74 63
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
6760 0 0
2
43514 0
0
5 4049~
219 607 714 0 2 22
0 14 76
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
5760 0 0
2
43514 0
0
5 4073~
219 990 687 0 4 22
0 77 11 76 75
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
3781 0 0
2
43514 0
0
5 4030~
219 853 644 0 3 22
0 15 72 77
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
8545 0 0
2
43514 0
0
14 Logic Display~
6 965 69 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9739 0 0
2
43514 0
0
14 Logic Display~
6 1013 70 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
388 0 0
2
43514 0
0
14 Logic Display~
6 1058 69 0 1 2
10 48
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4595 0 0
2
43514 0
0
14 Logic Display~
6 1100 67 0 1 2
10 66
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3173 0 0
2
43514 0
0
125
3 1 2 0 0 8320 0 14 13 0 0 7
2391 2971
2498 2971
2498 222
887 222
887 99
717 99
717 80
3 2 3 0 0 4224 0 15 14 0 0 4
2292 3010
2339 3010
2339 2980
2345 2980
3 1 4 0 0 8320 0 16 14 0 0 4
2320 2909
2336 2909
2336 2962
2345 2962
0 1 5 0 0 4096 0 0 15 14 0 5
1574 2600
1574 3045
1981 3045
1981 3001
2247 3001
0 2 6 0 0 8320 0 0 15 13 0 3
1682 2981
1682 3019
2247 3019
0 2 7 0 0 8320 0 0 16 11 0 3
1780 3181
1780 2918
2275 2918
3 1 8 0 0 8320 0 17 16 0 0 4
2253 2842
2269 2842
2269 2900
2275 2900
0 2 6 0 0 0 0 0 17 13 0 3
1816 2981
1816 2851
2204 2851
0 1 5 0 0 8320 0 0 17 14 0 3
1543 2600
1543 2833
2204 2833
3 1 9 0 0 8320 0 18 78 0 0 5
2119 3161
2142 3161
2142 140
965 140
965 87
3 2 7 0 0 0 0 21 18 0 0 4
1666 3181
2051 3181
2051 3170
2070 3170
3 1 10 0 0 8320 0 19 18 0 0 6
2061 3061
2082 3061
2082 3114
2039 3114
2039 3152
2070 3152
3 2 6 0 0 0 0 23 19 0 0 4
1630 2981
1963 2981
1963 3070
2012 3070
3 1 5 0 0 0 0 26 19 0 0 3
1444 2600
2012 2600
2012 3052
1 0 11 0 0 16512 0 20 0 0 122 8
1414 3164
1364 3164
1364 3322
1987 3322
1987 240
816 240
816 390
484 390
2 1 12 0 0 4224 0 20 21 0 0 4
1450 3164
1602 3164
1602 3172
1621 3172
3 2 13 0 0 8320 0 30 21 0 0 6
1465 2368
1894 2368
1894 3270
1580 3270
1580 3190
1621 3190
1 0 14 0 0 16512 0 24 0 0 120 8
1485 3012
1450 3012
1450 3103
1938 3103
1938 254
876 254
876 331
657 331
2 0 15 0 0 16512 0 25 0 0 125 6
1483 2962
1467 2962
1467 2772
1758 2772
1758 414
576 414
1 0 16 0 0 8192 0 22 0 0 22 3
1390 2936
1355 2936
1355 3030
2 1 17 0 0 4224 0 22 25 0 0 4
1426 2936
1460 2936
1460 2944
1483 2944
0 2 16 0 0 4096 0 0 24 32 0 3
1110 2527
1110 3030
1485 3030
3 2 18 0 0 4224 0 24 23 0 0 4
1530 3021
1572 3021
1572 2990
1584 2990
3 1 19 0 0 4224 0 25 23 0 0 4
1528 2953
1559 2953
1559 2972
1584 2972
1 2 20 0 0 8320 0 9 26 0 0 6
240 45
290 45
290 2925
1344 2925
1344 2609
1398 2609
4 1 21 0 0 4224 0 28 26 0 0 4
1276 2572
1345 2572
1345 2591
1398 2591
1 0 14 0 0 0 0 27 0 0 120 6
1022 2591
884 2591
884 2875
1721 2875
1721 353
657 353
2 0 11 0 0 0 0 28 0 0 122 6
1231 2572
1171 2572
1171 2679
1650 2679
1650 294
484 294
2 3 22 0 0 4224 0 27 28 0 0 3
1058 2591
1231 2591
1231 2581
3 1 23 0 0 8320 0 29 28 0 0 4
1192 2536
1210 2536
1210 2563
1231 2563
2 0 15 0 0 0 0 29 0 0 125 4
1143 2545
1081 2545
1081 269
576 269
1 1 16 0 0 8320 0 29 5 0 0 4
1143 2527
274 2527
274 111
243 111
3 2 24 0 0 8320 0 31 30 0 0 4
1382 2409
1411 2409
1411 2377
1419 2377
3 1 25 0 0 4224 0 32 30 0 0 4
1378 2344
1403 2344
1403 2359
1419 2359
0 2 26 0 0 12416 0 0 31 39 0 4
968 2138
958 2138
958 2418
1337 2418
0 1 27 0 0 8320 0 0 31 40 0 4
1029 1930
999 1930
999 2400
1337 2400
0 2 28 0 0 8320 0 0 32 42 0 3
940 2261
940 2353
1333 2353
3 1 29 0 0 8320 0 33 32 0 0 3
1270 2332
1270 2335
1333 2335
0 2 26 0 0 0 0 0 33 44 0 3
968 2105
968 2341
1221 2341
0 1 27 0 0 0 0 0 33 45 0 3
1029 1899
1029 2323
1221 2323
3 1 30 0 0 8320 0 34 79 0 0 5
1245 2072
1358 2072
1358 168
1013 168
1013 88
3 2 28 0 0 0 0 37 34 0 0 4
927 2261
1175 2261
1175 2081
1196 2081
3 1 31 0 0 12416 0 35 34 0 0 6
1199 1973
1228 1973
1228 2034
1161 2034
1161 2063
1196 2063
3 2 26 0 0 0 0 39 35 0 0 4
942 2105
1094 2105
1094 1982
1150 1982
3 1 27 0 0 0 0 42 35 0 0 4
1000 1899
1067 1899
1067 1964
1150 1964
1 0 11 0 0 0 0 36 0 0 122 4
712 2266
421 2266
421 357
484 357
2 2 32 0 0 4224 0 36 37 0 0 4
748 2266
839 2266
839 2270
882 2270
3 1 33 0 0 12416 0 46 37 0 0 6
1565 1554
1622 1554
1622 2202
830 2202
830 2252
882 2252
1 0 14 0 0 0 0 40 0 0 120 4
754 2141
458 2141
458 382
657 382
0 1 15 0 0 0 0 0 41 125 0 4
576 406
513 406
513 2048
752 2048
1 0 34 0 0 8192 0 38 0 0 53 3
649 2069
606 2069
606 2159
2 2 35 0 0 4224 0 38 41 0 0 4
685 2069
736 2069
736 2066
752 2066
0 2 34 0 0 4096 0 0 40 62 0 3
518 1834
518 2159
754 2159
3 2 36 0 0 4224 0 40 39 0 0 4
799 2150
865 2150
865 2114
896 2114
3 1 37 0 0 4224 0 41 39 0 0 4
797 2057
865 2057
865 2096
896 2096
1 2 38 0 0 16512 0 10 42 0 0 8
328 46
348 46
348 59
106 59
106 1963
915 1963
915 1908
954 1908
4 1 39 0 0 4224 0 44 42 0 0 4
854 1847
927 1847
927 1890
954 1890
0 1 14 0 0 0 0 0 43 120 0 6
657 475
608 475
608 1892
554 1892
554 1925
579 1925
2 3 40 0 0 4224 0 43 44 0 0 3
615 1925
809 1925
809 1856
0 2 11 0 0 0 0 0 44 77 0 5
254 431
254 1872
790 1872
790 1847
809 1847
3 1 41 0 0 4224 0 45 44 0 0 4
756 1825
796 1825
796 1838
809 1838
1 2 34 0 0 16512 0 6 45 0 0 6
325 112
343 112
343 145
21 145
21 1834
707 1834
0 1 15 0 0 0 0 0 45 125 0 4
576 480
40 480
40 1816
707 1816
2 3 42 0 0 8320 0 46 47 0 0 4
1519 1563
1506 1563
1506 1615
1471 1615
3 1 43 0 0 4224 0 48 46 0 0 4
1473 1511
1508 1511
1508 1545
1519 1545
0 2 44 0 0 8192 0 0 47 70 0 5
1126 1492
1126 1653
1414 1653
1414 1624
1426 1624
0 1 45 0 0 12416 0 0 47 71 0 4
1109 1353
1080 1353
1080 1606
1426 1606
0 2 46 0 0 4096 0 0 48 73 0 4
1185 1592
1417 1592
1417 1520
1428 1520
3 1 47 0 0 4224 0 49 48 0 0 4
1390 1483
1419 1483
1419 1502
1428 1502
0 2 44 0 0 8320 0 0 49 75 0 3
1044 1460
1044 1492
1341 1492
0 1 45 0 0 0 0 0 49 76 0 3
1109 1269
1109 1474
1341 1474
3 1 48 0 0 8320 0 50 80 0 0 5
1276 1421
1306 1421
1306 213
1058 213
1058 87
3 2 46 0 0 4224 0 53 50 0 0 4
914 1626
1185 1626
1185 1430
1227 1430
3 1 49 0 0 12416 0 51 50 0 0 6
1234 1340
1250 1340
1250 1379
1185 1379
1185 1412
1227 1412
3 2 44 0 0 0 0 55 51 0 0 4
1017 1460
1145 1460
1145 1349
1185 1349
3 1 45 0 0 0 0 58 51 0 0 4
1105 1269
1146 1269
1146 1331
1185 1331
1 0 11 0 0 0 0 52 0 0 122 4
638 1642
52 1642
52 431
484 431
2 2 50 0 0 4224 0 52 53 0 0 4
674 1642
855 1642
855 1635
869 1635
3 1 51 0 0 12416 0 62 53 0 0 6
1437 886
1492 886
1492 1565
811 1565
811 1617
869 1617
0 1 14 0 0 0 0 0 56 120 0 4
657 491
74 491
74 1495
880 1495
0 2 15 0 0 0 0 0 57 125 0 4
576 506
84 506
84 1432
878 1432
1 0 52 0 0 4096 0 54 0 0 84 3
673 1411
463 1411
463 1513
2 1 53 0 0 8320 0 54 57 0 0 3
709 1411
709 1414
878 1414
0 2 52 0 0 8320 0 0 56 94 0 4
207 441
96 441
96 1513
880 1513
3 2 54 0 0 8320 0 56 55 0 0 4
925 1504
944 1504
944 1469
971 1469
3 1 55 0 0 8320 0 57 55 0 0 4
923 1423
945 1423
945 1451
971 1451
1 2 56 0 0 16512 0 11 58 0 0 8
411 45
431 45
431 71
145 71
145 1304
1041 1304
1041 1278
1059 1278
4 1 57 0 0 8320 0 60 58 0 0 3
1009 1258
1009 1260
1059 1260
0 1 14 0 0 0 0 0 59 120 0 4
657 513
156 513
156 1279
727 1279
2 3 58 0 0 4224 0 59 60 0 0 4
763 1279
925 1279
925 1267
964 1267
0 2 11 0 0 0 0 0 60 122 0 4
484 530
166 530
166 1258
964 1258
3 1 59 0 0 4224 0 61 60 0 0 4
876 1227
924 1227
924 1249
964 1249
0 2 15 0 0 0 0 0 61 125 0 4
576 539
190 539
190 1236
827 1236
1 1 52 0 0 0 0 7 61 0 0 6
398 113
433 113
433 153
207 153
207 1218
827 1218
3 2 60 0 0 8320 0 63 62 0 0 4
1345 930
1366 930
1366 895
1391 895
3 1 61 0 0 4224 0 64 62 0 0 4
1335 847
1366 847
1366 877
1391 877
0 2 62 0 0 4224 0 0 63 101 0 4
1133 861
1261 861
1261 939
1300 939
0 1 63 0 0 12288 0 0 63 102 0 4
1139 772
1119 772
1119 921
1300 921
0 2 64 0 0 8320 0 0 64 104 0 5
1004 1036
1004 932
1272 932
1272 856
1290 856
3 1 65 0 0 4224 0 65 64 0 0 4
1213 814
1265 814
1265 838
1290 838
0 2 62 0 0 0 0 0 65 106 0 4
1094 892
1133 892
1133 823
1164 823
0 1 63 0 0 0 0 0 65 107 0 4
1101 748
1139 748
1139 805
1164 805
3 1 66 0 0 8320 0 66 81 0 0 5
1226 1045
1247 1045
1247 125
1100 125
1100 85
3 2 64 0 0 0 0 69 66 0 0 4
969 1036
1094 1036
1094 1054
1177 1054
3 1 67 0 0 8320 0 67 66 0 0 6
1168 974
1181 974
1181 1017
1151 1017
1151 1036
1177 1036
3 2 62 0 0 0 0 71 67 0 0 4
1086 872
1094 872
1094 983
1119 983
1 3 63 0 0 8320 0 67 74 0 0 4
1119 965
1101 965
1101 726
1079 726
1 2 68 0 0 20608 0 1 69 0 0 6
733 247
763 247
763 552
223 552
223 1045
924 1045
1 0 11 0 0 0 0 68 0 0 122 4
766 1027
242 1027
242 562
484 562
2 1 69 0 0 4224 0 68 69 0 0 2
802 1027
924 1027
2 0 14 0 0 0 0 73 0 0 120 4
916 844
269 844
269 572
657 572
0 2 15 0 0 0 0 0 72 125 0 4
576 584
285 584
285 924
920 924
3 2 70 0 0 4224 0 72 71 0 0 4
965 915
1012 915
1012 881
1040 881
3 1 71 0 0 4224 0 73 71 0 0 4
961 835
1010 835
1010 863
1040 863
0 1 72 0 0 8192 0 0 73 116 0 3
656 903
656 826
916 826
1 0 72 0 0 8320 0 70 0 0 124 4
751 903
352 903
352 157
537 157
2 1 73 0 0 8320 0 70 72 0 0 3
787 903
787 906
920 906
2 1 74 0 0 4224 0 74 12 0 0 6
1033 735
311 735
311 182
583 182
583 42
488 42
4 1 75 0 0 8320 0 76 74 0 0 4
1011 687
1027 687
1027 717
1033 717
1 1 14 0 0 0 0 4 75 0 0 6
638 253
657 253
657 593
386 593
386 714
592 714
2 3 76 0 0 4224 0 75 76 0 0 4
628 714
935 714
935 696
966 696
1 2 11 0 0 0 0 2 76 0 0 4
458 253
484 253
484 687
966 687
3 1 77 0 0 4224 0 77 76 0 0 4
886 644
934 644
934 678
966 678
1 2 72 0 0 0 0 8 77 0 0 6
490 109
537 109
537 205
406 205
406 653
837 653
1 1 15 0 0 0 0 3 77 0 0 4
558 255
576 255
576 635
837 635
26
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
656 108 757 132
666 116 746 132
10 Last Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2339 3016 2432 3040
2349 3024 2421 3040
9 CarryLast
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2077 3146 2114 3170
2087 3154 2103 3170
2 F3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1624 3166 1661 3190
1634 3174 1650 3190
2 Z3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1590 2967 1627 2991
1600 2975 1616 2991
2 Y3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1401 2583 1438 2607
1411 2591 1427 2607
2 X3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1423 2350 1460 2374
1433 2358 1449 2374
2 C2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1203 2053 1240 2077
1213 2061 1229 2077
2 F2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
888 2244 925 2268
898 2252 914 2268
2 Z2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
899 2088 936 2112
909 2096 925 2112
2 Y2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
955 1884 992 1908
965 1892 981 1908
2 X2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
588 1830 625 1854
598 1838 614 1854
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1522 1537 1559 1561
1532 1545 1548 1561
2 C1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1233 1405 1270 1429
1243 1413 1259 1429
2 F1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
870 1610 907 1634
880 1618 896 1634
2 Z1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
973 1442 1010 1466
983 1450 999 1466
2 Y1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1061 1253 1098 1277
1071 1261 1087 1277
2 X1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1393 869 1430 893
1403 877 1419 893
2 C0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1182 1030 1219 1054
1192 1038 1208 1054
2 F0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
928 1019 965 1043
938 1027 954 1043
2 Z0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1040 858 1077 882
1050 866 1066 882
2 Y0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1034 709 1071 733
1044 717 1060 733
2 X0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
943 13 980 37
953 21 969 37
2 F3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
993 10 1030 34
1003 18 1019 34
2 F2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1036 9 1073 33
1046 17 1062 33
2 F1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1081 7 1118 31
1091 15 1107 31
2 F0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
