CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 70 406 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 P5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4747 0 0
2
43548.4 0
0
13 Logic Switch~
5 73 343 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 P4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
972 0 0
2
43548.4 0
0
13 Logic Switch~
5 70 279 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 P3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3472 0 0
2
43548.4 0
0
13 Logic Switch~
5 72 238 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 P2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9998 0 0
2
43548.4 0
0
13 Logic Switch~
5 72 183 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 P1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3536 0 0
2
43548.4 0
0
13 Logic Switch~
5 72 131 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4597 0 0
2
43548.4 0
0
13 Logic Switch~
5 700 170 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 R
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3835 0 0
2
43548.4 0
0
13 Logic Switch~
5 71 75 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3670 0 0
2
43548.4 0
0
13 Logic Switch~
5 352 577 0 1 11
0 23
0
0 0 21360 0
2 0V
-14 -15 0 -7
5 clock
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5616 0 0
2
43548.4 0
0
9 2-In AND~
219 510 345 0 3 22
0 5 6 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
9323 0 0
2
43548.4 0
0
14 Logic Display~
6 949 148 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
317 0 0
2
43548.4 0
0
8 3-In OR~
219 352 411 0 4 22
0 2 8 7 6
0
0 0 624 0
4 4075
-14 -24 14 -16
4 Cout
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 5 0
1 U
3108 0 0
2
43548.4 0
0
9 2-In AND~
219 247 545 0 3 22
0 10 9 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
4299 0 0
2
43548.4 0
0
9 2-In AND~
219 246 468 0 3 22
0 11 10 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
9672 0 0
2
43548.4 0
0
9 2-In AND~
219 245 403 0 3 22
0 9 11 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7876 0 0
2
43548.4 0
0
8 4-In OR~
219 347 317 0 5 22
0 16 15 14 13 12
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
6369 0 0
2
43548.4 0
0
9 2-In AND~
219 254 346 0 3 22
0 11 17 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
9172 0 0
2
43548.4 0
0
8 3-In OR~
219 407 191 0 4 22
0 13 18 14 3
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 5 0
1 U
7100 0 0
2
43548.4 0
0
9 2-In AND~
219 325 238 0 3 22
0 11 19 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3820 0 0
2
43548.4 0
0
8 2-In OR~
219 198 228 0 3 22
0 17 20 19
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7678 0 0
2
43548.4 0
0
9 2-In AND~
219 292 77 0 3 22
0 21 5 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
961 0 0
2
43548.4 0
0
9 2-In XOR~
219 201 105 0 3 22
0 11 10 21
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3178 0 0
2
43548.4 0
0
14 Logic Display~
6 1024 77 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3409 0 0
2
43548.4 0
0
7 Pulser~
4 440 506 0 11 12
0 23 25 24 26 0 0 5 5 -1
7 1
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3951 0 0
2
43548.4 0
0
6 JK RN~
219 761 95 0 6 22
0 3 24 12 22 27 9
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
8885 0 0
2
43548.4 0
0
35
3 1 2 0 0 8320 0 15 12 0 0 3
266 403
266 402
339 402
4 1 3 0 0 12416 0 18 25 0 0 4
440 191
563 191
563 78
737 78
3 1 4 0 0 4224 0 10 11 0 0 3
531 345
949 345
949 166
0 1 5 0 0 8320 0 0 10 28 0 4
251 111
461 111
461 336
486 336
4 2 6 0 0 4224 0 12 10 0 0 4
385 411
480 411
480 354
486 354
3 3 7 0 0 4224 0 13 12 0 0 3
268 545
268 420
339 420
3 2 8 0 0 8320 0 14 12 0 0 4
267 468
289 468
289 411
340 411
0 2 9 0 0 4096 0 0 13 12 0 3
200 391
200 554
223 554
0 1 10 0 0 8192 0 0 13 10 0 3
107 477
107 536
223 536
0 2 10 0 0 4224 0 0 14 30 0 3
107 131
107 477
222 477
0 1 11 0 0 8192 0 0 14 13 0 3
114 412
114 459
222 459
0 1 9 0 0 8320 0 0 15 33 0 5
886 95
886 370
200 370
200 394
221 394
0 2 11 0 0 0 0 0 15 19 0 3
114 335
114 412
221 412
5 3 12 0 0 4224 0 16 25 0 0 4
380 317
632 317
632 96
737 96
0 4 13 0 0 8320 0 0 16 24 0 4
377 137
287 137
287 331
330 331
0 3 14 0 0 8192 0 0 16 22 0 3
243 279
243 322
330 322
1 2 15 0 0 12416 0 4 16 0 0 6
84 238
132 238
132 265
295 265
295 313
330 313
3 1 16 0 0 8320 0 17 16 0 0 3
275 346
275 304
330 304
0 1 11 0 0 4224 0 0 17 31 0 3
114 75
114 337
230 337
0 1 11 0 0 0 0 0 19 31 0 5
163 94
163 191
280 191
280 229
301 229
0 2 17 0 0 12288 0 0 17 27 0 4
144 343
155 343
155 355
230 355
1 3 14 0 0 4224 0 3 18 0 0 4
82 279
380 279
380 200
394 200
3 2 18 0 0 8320 0 19 18 0 0 4
346 238
361 238
361 191
395 191
3 1 13 0 0 0 0 21 18 0 0 4
313 77
377 77
377 182
394 182
3 2 19 0 0 12416 0 20 19 0 0 4
231 228
262 228
262 247
301 247
1 2 20 0 0 8320 0 1 20 0 0 4
82 406
165 406
165 237
185 237
1 1 17 0 0 8320 0 2 20 0 0 4
85 343
147 343
147 219
185 219
1 2 5 0 0 128 0 5 21 0 0 4
84 183
251 183
251 86
268 86
3 1 21 0 0 8320 0 22 21 0 0 4
234 105
243 105
243 68
268 68
1 2 10 0 0 0 0 6 22 0 0 4
84 131
137 131
137 114
185 114
1 1 11 0 0 0 0 8 22 0 0 4
83 75
163 75
163 96
185 96
1 4 22 0 0 4224 0 7 25 0 0 3
712 170
761 170
761 126
6 1 9 0 0 128 0 25 23 0 0 4
785 78
798 78
798 95
1024 95
1 1 23 0 0 8320 0 24 9 0 0 3
416 497
364 497
364 577
3 2 24 0 0 8320 0 24 25 0 0 4
464 497
588 497
588 87
730 87
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
