CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
3 100 1 2 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
41
13 Logic Switch~
5 662 331 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3171 0 0
2
43537 0
0
13 Logic Switch~
5 470 331 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4139 0 0
2
43537 0
0
13 Logic Switch~
5 561 334 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6435 0 0
2
43537 0
0
13 Logic Switch~
5 189 201 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5283 0 0
2
43537 0
0
13 Logic Switch~
5 334 195 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6874 0 0
2
43537 0
0
13 Logic Switch~
5 188 111 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5305 0 0
2
43537 0
0
13 Logic Switch~
5 337 107 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
34 0 0
2
43537 0
0
5 4071~
219 1205 1231 0 3 22
0 3 4 2
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U10B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 10 0
1 U
969 0 0
2
43537 0
0
5 4081~
219 1080 1280 0 3 22
0 6 5 4
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 7 0
1 U
8402 0 0
2
43537 0
0
5 4081~
219 906 1400 0 3 22
0 8 7 3
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 7 0
1 U
3751 0 0
2
43537 0
0
5 4030~
219 1121 1464 0 3 22
0 6 5 9
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U6D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 6 0
1 U
4292 0 0
2
43537 0
0
5 4030~
219 992 1368 0 3 22
0 8 7 6
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U6C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 6 0
1 U
6118 0 0
2
43537 0
0
5 4071~
219 874 1581 0 3 22
0 11 10 7
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 10 0
1 U
34 0 0
2
43537 0
0
5 4049~
219 445 1708 0 2 22
0 12 13
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 8 0
1 U
6357 0 0
2
43537 0
0
5 4073~
219 586 1689 0 4 22
0 15 14 13 10
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 9 0
1 U
319 0 0
2
43537 0
0
5 4049~
219 624 1521 0 2 22
0 15 16
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 8 0
1 U
3976 0 0
2
43537 0
0
5 4081~
219 750 1513 0 3 22
0 17 16 11
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
7634 0 0
2
43537 0
0
5 4071~
219 797 1267 0 3 22
0 19 18 8
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
523 0 0
2
43537 0
0
5 4049~
219 475 1359 0 2 22
0 12 20
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
6748 0 0
2
43537 0
0
5 4049~
219 560 1319 0 2 22
0 21 22
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
6901 0 0
2
43537 0
0
5 4073~
219 670 1331 0 4 22
0 22 14 20 18
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 2 0
1 U
842 0 0
2
43537 0
0
5 4081~
219 670 1219 0 3 22
0 12 21 19
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
3277 0 0
2
43537 0
0
5 4071~
219 1042 737 0 3 22
0 24 23 5
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
4212 0 0
2
43537 0
0
5 4081~
219 1023 794 0 3 22
0 25 26 23
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
4720 0 0
2
43537 0
0
5 4081~
219 997 713 0 3 22
0 28 27 24
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
5551 0 0
2
43537 0
0
5 4030~
219 1000 1036 0 3 22
0 26 25 29
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
6986 0 0
2
43537 0
0
5 4030~
219 919 993 0 3 22
0 28 27 26
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
8745 0 0
2
43537 0
0
5 4071~
219 796 901 0 3 22
0 31 30 27
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
9592 0 0
2
43537 0
0
5 4049~
219 468 965 0 2 22
0 12 32
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
8748 0 0
2
43537 0
0
5 4073~
219 698 951 0 4 22
0 33 14 32 30
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
7168 0 0
2
43537 0
0
5 4049~
219 503 870 0 2 22
0 33 34
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
631 0 0
2
43537 0
0
5 4081~
219 699 857 0 3 22
0 17 34 31
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
9466 0 0
2
43537 0
0
10 2-In XNOR~
219 567 826 0 3 22
0 12 14 17
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U5A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
3266 0 0
2
43537 0
0
5 4071~
219 599 534 0 3 22
0 36 35 28
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
7693 0 0
2
43537 0
0
5 4049~
219 348 630 0 2 22
0 12 37
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
3723 0 0
2
43537 0
0
5 4049~
219 371 584 0 2 22
0 38 39
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
3440 0 0
2
43537 0
0
5 4073~
219 479 593 0 4 22
0 39 14 37 35
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
6263 0 0
2
43537 0
0
5 4081~
219 474 473 0 3 22
0 12 38 36
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
4900 0 0
2
43537 0
0
14 Logic Display~
6 655 73 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8783 0 0
2
43537 0
0
14 Logic Display~
6 895 67 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3221 0 0
2
43537 0
0
14 Logic Display~
6 981 65 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3215 0 0
2
43537 0
0
61
3 1 2 0 0 8320 0 8 39 0 0 5
1238 1231
1309 1231
1309 126
655 126
655 91
3 1 3 0 0 4224 0 10 8 0 0 4
927 1400
1167 1400
1167 1222
1192 1222
3 2 4 0 0 4224 0 9 8 0 0 4
1101 1280
1164 1280
1164 1240
1192 1240
0 2 5 0 0 8192 0 0 9 9 0 4
1121 1155
1001 1155
1001 1289
1056 1289
0 1 6 0 0 4224 0 0 9 10 0 3
1041 1368
1041 1271
1056 1271
0 2 7 0 0 4096 0 0 10 11 0 5
912 1581
912 1459
853 1459
853 1409
882 1409
0 1 8 0 0 4224 0 0 10 12 0 3
845 1267
845 1391
882 1391
3 1 9 0 0 8320 0 11 40 0 0 5
1154 1464
1280 1464
1280 161
895 161
895 85
3 2 5 0 0 8320 0 23 11 0 0 6
1075 737
1121 737
1121 1415
1046 1415
1046 1473
1105 1473
3 1 6 0 0 0 0 12 11 0 0 4
1025 1368
1075 1368
1075 1455
1105 1455
3 2 7 0 0 8320 0 13 12 0 0 4
907 1581
964 1581
964 1377
976 1377
3 1 8 0 0 0 0 18 12 0 0 4
830 1267
932 1267
932 1359
976 1359
4 2 10 0 0 4224 0 15 13 0 0 4
607 1689
815 1689
815 1590
861 1590
3 1 11 0 0 8320 0 17 13 0 0 4
771 1513
814 1513
814 1572
861 1572
1 0 12 0 0 8320 0 14 0 0 61 4
430 1708
328 1708
328 388
502 388
2 3 13 0 0 4224 0 14 15 0 0 4
466 1708
532 1708
532 1698
562 1698
0 2 14 0 0 4224 0 0 15 57 0 5
559 417
559 1643
400 1643
400 1689
562 1689
0 1 15 0 0 4096 0 0 15 19 0 3
442 1521
442 1680
562 1680
1 1 15 0 0 8320 0 16 4 0 0 6
609 1521
78 1521
78 241
218 241
218 201
201 201
2 2 16 0 0 8320 0 16 17 0 0 3
645 1521
645 1522
726 1522
0 1 17 0 0 4224 0 0 17 50 0 3
613 826
613 1504
726 1504
4 2 18 0 0 4224 0 21 18 0 0 4
691 1331
759 1331
759 1276
784 1276
3 1 19 0 0 4224 0 22 18 0 0 4
691 1219
752 1219
752 1258
784 1258
1 0 12 0 0 0 0 19 0 0 61 4
460 1359
296 1359
296 343
502 343
2 3 20 0 0 4224 0 19 21 0 0 4
496 1359
631 1359
631 1340
646 1340
0 2 14 0 0 0 0 0 21 57 0 4
597 361
212 361
212 1331
646 1331
1 0 21 0 0 4096 0 20 0 0 29 3
545 1319
352 1319
352 1228
2 1 22 0 0 8320 0 20 21 0 0 3
581 1319
581 1322
646 1322
1 2 21 0 0 8320 0 6 22 0 0 4
200 111
282 111
282 1228
646 1228
0 1 12 0 0 0 0 0 22 44 0 3
430 350
430 1210
646 1210
2 3 23 0 0 12416 0 23 24 0 0 6
1029 746
1015 746
1015 761
1067 761
1067 794
1044 794
3 1 24 0 0 8320 0 25 23 0 0 4
1018 713
1025 713
1025 728
1029 728
0 1 25 0 0 4096 0 0 24 38 0 3
851 331
851 785
999 785
0 2 26 0 0 8320 0 0 24 39 0 4
975 1000
987 1000
987 803
999 803
0 2 27 0 0 4224 0 0 25 40 0 3
844 901
844 722
973 722
0 1 28 0 0 8192 0 0 25 41 0 3
792 534
792 704
973 704
3 1 29 0 0 8320 0 26 41 0 0 5
1033 1036
1094 1036
1094 102
981 102
981 83
2 1 25 0 0 8320 0 26 1 0 0 4
984 1045
956 1045
956 331
674 331
3 1 26 0 0 0 0 27 26 0 0 4
952 993
975 993
975 1027
984 1027
3 2 27 0 0 0 0 28 27 0 0 4
829 901
855 901
855 1002
903 1002
3 1 28 0 0 8320 0 34 27 0 0 4
632 534
897 534
897 984
903 984
4 2 30 0 0 4224 0 30 28 0 0 4
719 951
768 951
768 910
783 910
3 1 31 0 0 8320 0 32 28 0 0 4
720 857
748 857
748 892
783 892
1 0 12 0 0 0 0 29 0 0 61 4
453 965
27 965
27 350
502 350
2 3 32 0 0 4224 0 29 30 0 0 4
489 965
650 965
650 960
674 960
0 2 14 0 0 0 0 0 30 57 0 4
597 377
49 377
49 951
674 951
0 1 33 0 0 8192 0 0 30 48 0 3
279 870
279 942
674 942
1 1 33 0 0 8320 0 31 5 0 0 6
488 870
88 870
88 335
364 335
364 195
346 195
2 2 34 0 0 4224 0 31 32 0 0 4
524 870
667 870
667 866
675 866
3 1 17 0 0 0 0 33 32 0 0 4
606 826
639 826
639 848
675 848
0 2 14 0 0 0 0 0 33 57 0 4
597 396
117 396
117 835
551 835
0 1 12 0 0 0 0 0 33 55 0 4
250 432
148 432
148 817
551 817
4 2 35 0 0 8320 0 37 34 0 0 4
500 593
541 593
541 543
586 543
3 1 36 0 0 8320 0 38 34 0 0 4
495 473
541 473
541 525
586 525
1 0 12 0 0 0 0 35 0 0 61 4
333 630
250 630
250 369
502 369
2 3 37 0 0 4224 0 35 37 0 0 4
369 630
430 630
430 602
455 602
1 2 14 0 0 0 0 3 37 0 0 8
573 334
597 334
597 417
321 417
321 607
407 607
407 593
455 593
1 0 38 0 0 4096 0 36 0 0 60 3
356 584
356 443
398 443
2 1 39 0 0 4224 0 36 37 0 0 2
392 584
455 584
1 2 38 0 0 8320 0 7 38 0 0 4
349 107
398 107
398 482
450 482
1 1 12 0 0 0 0 2 38 0 0 6
482 331
502 331
502 406
412 406
412 464
450 464
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1192 1213 1229 1237
1202 1221 1218 1237
2 C1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1112 1446 1149 1470
1122 1454 1138 1470
2 F1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
863 1566 900 1590
873 1574 889 1590
2 Y1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
786 1251 823 1275
796 1259 812 1275
2 X1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1032 718 1069 742
1042 726 1058 742
2 C0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
991 1021 1028 1045
1001 1029 1017 1045
2 F0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
784 883 821 907
794 891 810 907
2 Y0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
587 517 624 541
597 525 613 541
2 X0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
548 20 649 44
558 28 638 44
10 Carry Last
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
873 4 910 28
883 12 899 28
2 F1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
962 4 999 28
972 12 988 28
2 F0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
