CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
3 100 1 2 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
44
13 Logic Switch~
5 581 266 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4797 0 0
2
43534.9 0
0
13 Logic Switch~
5 369 271 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4681 0 0
2
43534.9 0
0
13 Logic Switch~
5 474 274 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9730 0 0
2
43534.9 0
0
13 Logic Switch~
5 149 161 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9874 0 0
2
43534.9 0
0
13 Logic Switch~
5 233 163 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
364 0 0
2
43534.9 0
0
13 Logic Switch~
5 148 88 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3656 0 0
2
43534.9 0
0
13 Logic Switch~
5 234 84 0 1 11
0 38
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3131 0 0
2
43534.9 0
0
5 4071~
219 1162 1488 0 3 22
0 5 4 3
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 7 0
1 U
6772 0 0
2
43534.9 0
0
5 4081~
219 1069 1476 0 3 22
0 7 6 5
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U8D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 8 0
1 U
9557 0 0
2
43534.9 0
0
5 4081~
219 1107 1542 0 3 22
0 8 2 4
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U8C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 8 0
1 U
5789 0 0
2
43534.9 0
0
14 Logic Display~
6 572 57 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7328 0 0
2
43534.9 0
0
5 4030~
219 1065 1419 0 3 22
0 8 2 9
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U5D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
4799 0 0
2
43534.9 0
0
5 4030~
219 942 1340 0 3 22
0 7 6 8
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U5C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
9196 0 0
2
43534.9 0
0
5 4071~
219 884 1527 0 3 22
0 11 10 6
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 7 0
1 U
3857 0 0
2
43534.9 0
0
5 4049~
219 560 1642 0 2 22
0 12 13
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 6 0
1 U
7125 0 0
2
43534.9 0
0
5 4049~
219 592 1610 0 2 22
0 15 16
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 6 0
1 U
3641 0 0
2
43534.9 0
0
5 4073~
219 695 1620 0 4 22
0 16 14 13 10
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 9 0
1 U
9821 0 0
2
43534.9 0
0
5 4081~
219 774 1452 0 3 22
0 12 15 11
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 8 0
1 U
3187 0 0
2
43534.9 0
0
5 4071~
219 726 1222 0 3 22
0 18 17 7
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
762 0 0
2
43534.9 0
0
5 4081~
219 602 1305 0 3 22
0 20 19 17
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 8 0
1 U
39 0 0
2
43534.9 0
0
5 4049~
219 368 1250 0 2 22
0 12 21
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 6 0
1 U
9450 0 0
2
43534.9 0
0
5 4071~
219 483 1255 0 3 22
0 21 14 20
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
3236 0 0
2
43534.9 0
0
5 4049~
219 369 1155 0 2 22
0 14 22
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 6 0
1 U
3321 0 0
2
43534.9 0
0
5 4049~
219 410 1128 0 2 22
0 19 23
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 2 0
1 U
8879 0 0
2
43534.9 0
0
5 4073~
219 495 1136 0 4 22
0 23 22 12 18
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 1 0
1 U
5433 0 0
2
43534.9 0
0
5 4071~
219 1106 888 0 3 22
0 25 24 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
3679 0 0
2
43534.9 0
0
5 4081~
219 1013 764 0 3 22
0 27 26 25
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
9342 0 0
2
43534.9 0
0
5 4081~
219 1012 1048 0 3 22
0 29 28 24
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
3623 0 0
2
43534.9 0
0
5 4030~
219 991 917 0 3 22
0 29 28 30
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U5B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
3722 0 0
2
43534.9 0
0
5 4030~
219 909 888 0 3 22
0 27 26 29
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U5A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
8993 0 0
2
43534.9 0
0
5 4071~
219 792 698 0 3 22
0 32 31 26
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
3723 0 0
2
43534.9 0
0
5 4049~
219 536 762 0 2 22
0 12 33
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 2 0
1 U
6244 0 0
2
43534.9 0
0
5 4049~
219 588 731 0 2 22
0 34 35
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 2 0
1 U
6421 0 0
2
43534.9 0
0
5 4073~
219 668 742 0 4 22
0 35 14 33 31
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 1 0
1 U
7743 0 0
2
43534.9 0
0
5 4081~
219 670 670 0 3 22
0 12 34 32
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
9840 0 0
2
43534.9 0
0
5 4071~
219 842 493 0 3 22
0 37 36 27
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
6910 0 0
2
43534.9 0
0
5 4081~
219 824 592 0 3 22
0 39 38 36
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
449 0 0
2
43534.9 0
0
5 4049~
219 587 567 0 2 22
0 12 40
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 2 0
1 U
8761 0 0
2
43534.9 0
0
5 4071~
219 688 555 0 3 22
0 14 40 39
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
6748 0 0
2
43534.9 0
0
5 4049~
219 561 469 0 2 22
0 14 41
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 2 0
1 U
7393 0 0
2
43534.9 0
0
5 4049~
219 562 439 0 2 22
0 38 42
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 2 0
1 U
7699 0 0
2
43534.9 0
0
5 4073~
219 701 451 0 4 22
0 42 41 12 37
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 1 0
1 U
6638 0 0
2
43534.9 0
0
14 Logic Display~
6 858 54 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4595 0 0
2
43534.9 0
0
14 Logic Display~
6 924 51 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9395 0 0
2
43534.9 0
0
65
0 2 2 0 0 16512 0 0 10 9 0 8
1153 964
1127 964
1127 1022
1389 1022
1389 1591
1059 1591
1059 1551
1083 1551
3 1 3 0 0 8320 0 8 11 0 0 5
1195 1488
1281 1488
1281 204
572 204
572 75
3 2 4 0 0 8320 0 10 8 0 0 4
1128 1542
1142 1542
1142 1497
1149 1497
3 1 5 0 0 4224 0 9 8 0 0 4
1090 1476
1136 1476
1136 1479
1149 1479
0 2 6 0 0 8192 0 0 9 11 0 3
952 1484
952 1485
1045 1485
0 1 7 0 0 8320 0 0 9 12 0 3
864 1331
864 1467
1045 1467
0 1 8 0 0 4224 0 0 10 10 0 3
978 1340
978 1533
1083 1533
3 1 9 0 0 8320 0 12 43 0 0 5
1098 1419
1166 1419
1166 159
858 159
858 72
3 2 2 0 0 128 0 26 12 0 0 6
1139 888
1153 888
1153 1360
997 1360
997 1428
1049 1428
3 1 8 0 0 128 0 13 12 0 0 6
975 1340
1047 1340
1047 1378
1033 1378
1033 1410
1049 1410
3 2 6 0 0 8320 0 14 13 0 0 6
917 1527
952 1527
952 1379
895 1379
895 1349
926 1349
3 1 7 0 0 128 0 19 13 0 0 4
759 1222
847 1222
847 1331
926 1331
4 2 10 0 0 4224 0 17 14 0 0 4
716 1620
852 1620
852 1536
871 1536
3 1 11 0 0 8320 0 18 14 0 0 4
795 1452
828 1452
828 1518
871 1518
1 0 12 0 0 16384 0 15 0 0 61 8
545 1642
363 1642
363 1349
299 1349
299 278
348 278
348 288
416 288
2 3 13 0 0 4224 0 15 17 0 0 4
581 1642
664 1642
664 1629
671 1629
0 2 14 0 0 8320 0 0 17 62 0 4
496 377
174 377
174 1620
671 1620
1 0 15 0 0 8192 0 16 0 0 20 3
577 1610
488 1610
488 1461
2 1 16 0 0 8320 0 16 17 0 0 3
613 1610
613 1611
671 1611
1 2 15 0 0 16512 0 4 18 0 0 6
161 161
181 161
181 181
24 181
24 1461
750 1461
0 1 12 0 0 8320 0 0 18 61 0 4
416 364
67 364
67 1443
750 1443
2 3 17 0 0 8320 0 19 20 0 0 4
713 1231
653 1231
653 1305
623 1305
4 1 18 0 0 4224 0 25 19 0 0 4
516 1136
690 1136
690 1213
713 1213
2 0 19 0 0 8320 0 20 0 0 32 4
578 1314
115 1314
115 109
200 109
3 1 20 0 0 8320 0 22 20 0 0 4
516 1255
553 1255
553 1296
578 1296
0 2 14 0 0 0 0 0 22 62 0 6
496 308
205 308
205 1267
461 1267
461 1264
470 1264
1 0 12 0 0 0 0 21 0 0 61 4
353 1250
266 1250
266 331
416 331
2 1 21 0 0 4224 0 21 22 0 0 4
389 1250
460 1250
460 1246
470 1246
0 3 12 0 0 0 0 0 25 61 0 6
416 386
221 386
221 1188
462 1188
462 1145
471 1145
1 0 14 0 0 0 0 23 0 0 62 6
354 1155
305 1155
305 503
324 503
324 409
496 409
2 2 22 0 0 4224 0 23 25 0 0 4
390 1155
445 1155
445 1136
471 1136
1 1 19 0 0 0 0 24 6 0 0 6
395 1128
158 1128
158 210
200 210
200 88
160 88
2 1 23 0 0 8320 0 24 25 0 0 3
431 1128
431 1127
471 1127
3 2 24 0 0 8320 0 28 26 0 0 4
1033 1048
1087 1048
1087 897
1093 897
3 1 25 0 0 8320 0 27 26 0 0 4
1034 764
1086 764
1086 879
1093 879
0 2 26 0 0 4096 0 0 27 43 0 2
844 773
989 773
0 1 27 0 0 4096 0 0 27 44 0 4
899 736
979 736
979 755
989 755
0 2 28 0 0 4096 0 0 28 41 0 3
970 926
970 1057
988 1057
0 1 29 0 0 4224 0 0 28 42 0 3
955 888
955 1039
988 1039
3 1 30 0 0 8320 0 29 44 0 0 5
1024 917
1073 917
1073 95
924 95
924 69
1 2 28 0 0 8320 0 1 29 0 0 6
593 266
937 266
937 848
945 848
945 926
975 926
3 1 29 0 0 0 0 30 29 0 0 4
942 888
964 888
964 908
975 908
3 2 26 0 0 8320 0 31 30 0 0 4
825 698
844 698
844 897
893 897
3 1 27 0 0 8320 0 36 30 0 0 6
875 493
899 493
899 847
853 847
853 879
893 879
4 2 31 0 0 4224 0 34 31 0 0 4
689 742
772 742
772 707
779 707
3 1 32 0 0 4224 0 35 31 0 0 4
691 670
762 670
762 689
779 689
1 0 12 0 0 0 0 32 0 0 58 3
521 762
466 762
466 567
2 3 33 0 0 4224 0 32 34 0 0 4
557 762
628 762
628 751
644 751
0 2 14 0 0 0 0 0 34 62 0 3
524 469
524 742
644 742
1 0 34 0 0 4096 0 33 0 0 52 3
573 731
516 731
516 679
2 1 35 0 0 8320 0 33 34 0 0 3
609 731
609 733
644 733
1 2 34 0 0 8320 0 5 35 0 0 4
245 163
284 163
284 679
646 679
0 1 12 0 0 0 0 0 35 58 0 3
499 567
499 661
646 661
3 2 36 0 0 8320 0 37 36 0 0 6
845 592
860 592
860 528
805 528
805 502
829 502
4 1 37 0 0 4224 0 42 36 0 0 4
722 451
799 451
799 484
829 484
0 2 38 0 0 8320 0 0 37 64 0 3
347 439
347 601
800 601
3 1 39 0 0 4224 0 39 37 0 0 4
721 555
778 555
778 583
800 583
1 0 12 0 0 0 0 38 0 0 61 3
572 567
448 567
448 488
2 2 40 0 0 4224 0 38 39 0 0 4
608 567
655 567
655 564
675 564
0 1 14 0 0 0 0 0 39 62 0 3
540 469
540 546
675 546
1 3 12 0 0 0 0 2 42 0 0 6
381 271
416 271
416 488
655 488
655 460
677 460
1 1 14 0 0 0 0 40 3 0 0 4
546 469
496 469
496 274
486 274
2 2 41 0 0 12416 0 40 42 0 0 4
582 469
627 469
627 451
677 451
1 1 38 0 0 0 0 41 7 0 0 4
547 439
303 439
303 84
246 84
2 1 42 0 0 8320 0 41 42 0 0 3
583 439
583 442
677 442
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
464 39 565 63
474 47 554 63
10 Carry Last
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1053 1404 1090 1428
1063 1412 1079 1428
2 F1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
873 1513 910 1537
883 1521 899 1537
2 Y1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
715 1204 752 1228
725 1212 741 1228
2 X1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1095 871 1132 895
1105 879 1121 895
2 C0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
875 920 976 944
885 928 965 944
10 Cin Direct
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
980 899 1017 923
990 907 1006 923
2 F0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
784 682 821 706
794 690 810 706
2 Y0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
832 476 869 500
842 484 858 500
2 X0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
838 0 875 24
848 8 864 24
2 F1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
905 0 942 24
915 8 931 24
2 F0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
