CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9961490 0
0
6 Title:
5 Name:
0
0
0
64
5 4030~
219 1214 3369 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
4 U13A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 13 0
1 U
5616 0 0
2
43514 15
0
5 4071~
219 1606 3215 0 1 22
0 0
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U8D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 8 0
1 U
9323 0 0
2
43514 14
0
5 4081~
219 1520 3240 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
4 U12C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 12 0
1 U
317 0 0
2
43514 13
0
5 4081~
219 1519 3194 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
4 U12B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 12 0
1 U
3108 0 0
2
43514 12
0
5 4030~
219 1370 3177 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
4 U10D
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 10 0
1 U
4299 0 0
2
43514 11
0
5 4030~
219 1632 2729 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
4 U10C
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 10 0
1 U
9672 0 0
2
43514 10
0
5 4030~
219 1611 2602 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
4 U10B
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 10 0
1 U
7876 0 0
2
43514 9
0
5 4049~
219 773 2905 0 1 22
0 0
0
0 0 608 0
4 4049
-7 -24 21 -16
4 U11C
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 11 0
1 U
6369 0 0
2
43514 8
0
5 4081~
219 925 2916 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
4 U12A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 12 0
1 U
9172 0 0
2
43514 7
0
5 4049~
219 726 2669 0 1 22
0 0
0
0 0 608 0
4 4049
-7 -24 21 -16
4 U11B
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 11 0
1 U
7100 0 0
2
43514 6
0
5 4071~
219 1057 2726 0 1 22
0 0
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 8 0
1 U
3820 0 0
2
43514 5
0
5 4081~
219 951 2761 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 9 0
1 U
7678 0 0
2
43514 4
0
5 4081~
219 950 2686 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 9 0
1 U
961 0 0
2
43514 3
0
5 4049~
219 912 2543 0 1 22
0 0
0
0 0 608 0
4 4049
-7 -24 21 -16
4 U11A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 11 0
1 U
3178 0 0
2
43514 2
0
5 4073~
219 1132 2514 0 1 22
0 0
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 2 0
1 U
3409 0 0
2
43514 1
0
5 4030~
219 1051 2434 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
4 U10A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 10 0
1 U
3951 0 0
2
43514 0
0
5 4071~
219 1363 2207 0 1 22
0 0
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 8 0
1 U
8885 0 0
2
43514 47
0
5 4081~
219 1248 2245 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 9 0
1 U
3780 0 0
2
43514 46
0
5 4081~
219 1246 2175 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 9 0
1 U
9265 0 0
2
43514 45
0
5 4030~
219 1106 2152 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U7D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 7 0
1 U
9442 0 0
2
43514 44
0
5 4030~
219 1248 1944 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U7C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 7 0
1 U
9424 0 0
2
43514 43
0
5 4030~
219 1201 1818 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U7B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
9968 0 0
2
43514 42
0
5 4049~
219 880 1925 0 1 22
0 0
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U3F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
9281 0 0
2
43514 41
0
5 4081~
219 1011 1928 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 6 0
1 U
8464 0 0
2
43514 40
0
5 4071~
219 1088 1730 0 1 22
0 0
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 8 0
1 U
7168 0 0
2
43514 39
0
5 4049~
219 781 1679 0 1 22
0 0
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U3E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
3171 0 0
2
43514 38
0
5 4081~
219 991 1776 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 6 0
1 U
4139 0 0
2
43514 37
0
5 4081~
219 989 1697 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
6435 0 0
2
43514 36
0
5 4071~
219 996 1600 0 1 22
0 0
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
5283 0 0
2
43514 35
0
5 4049~
219 649 1487 0 1 22
0 0
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
6874 0 0
2
43514 34
0
5 4073~
219 887 1442 0 1 22
0 0
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
5305 0 0
2
43514 33
0
5 4030~
219 749 1376 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U7A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
34 0 0
2
43514 32
0
5 4071~
219 1076 1097 0 1 22
0 0
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
969 0 0
2
43514 31
0
5 4081~
219 1012 1134 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
8402 0 0
2
43514 30
0
5 4081~
219 1007 1066 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
3751 0 0
2
43514 29
0
5 4030~
219 953 976 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
4292 0 0
2
43514 28
0
5 4030~
219 1040 752 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
6118 0 0
2
43514 27
0
5 4030~
219 1004 647 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
34 0 0
2
43514 26
0
14 Logic Display~
6 1014 63 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6357 0 0
2
43514 25
0
14 Logic Display~
6 1056 62 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
319 0 0
2
43514 24
0
14 Logic Display~
6 1094 62 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3976 0 0
2
43514 23
0
14 Logic Display~
6 1134 62 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7634 0 0
2
43514 22
0
5 4049~
219 794 852 0 1 22
0 0
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
523 0 0
2
43514 21
0
5 4081~
219 913 837 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
6748 0 0
2
43514 20
0
5 4071~
219 909 699 0 1 22
0 0
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
6901 0 0
2
43514 19
0
5 4049~
219 570 649 0 1 22
0 0
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
842 0 0
2
43514 18
0
5 4081~
219 719 744 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
3277 0 0
2
43514 17
0
5 4081~
219 723 655 0 1 22
0 0
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
4212 0 0
2
43514 16
0
5 4071~
219 911 593 0 1 22
0 0
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
4720 0 0
2
43514 15
0
5 4049~
219 618 603 0 1 22
0 0
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
5551 0 0
2
43514 14
0
5 4073~
219 823 579 0 1 22
0 0
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
6986 0 0
2
43514 13
0
5 4030~
219 692 530 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
8745 0 0
2
43514 12
0
13 Logic Switch~
5 706 389 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9592 0 0
2
43514 11
0
13 Logic Switch~
5 423 399 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 S2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8748 0 0
2
43514 10
0
13 Logic Switch~
5 523 402 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7168 0 0
2
43514 9
0
13 Logic Switch~
5 602 403 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
631 0 0
2
43514 8
0
13 Logic Switch~
5 151 184 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9466 0 0
2
43514 7
0
13 Logic Switch~
5 266 185 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3266 0 0
2
43514 6
0
13 Logic Switch~
5 375 187 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7693 0 0
2
43514 5
0
13 Logic Switch~
5 486 185 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3723 0 0
2
43514 4
0
13 Logic Switch~
5 146 75 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3440 0 0
2
43514 3
0
13 Logic Switch~
5 264 79 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6263 0 0
2
43514 2
0
13 Logic Switch~
5 380 79 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4900 0 0
2
43514 1
0
13 Logic Switch~
5 482 77 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8783 0 0
2
43514 0
0
91
3 2 0 0 0 16 0 3 2 0 0 4
1541 3240
1568 3240
1568 3224
1593 3224
3 1 0 0 0 16 0 4 2 0 0 4
1540 3194
1567 3194
1567 3206
1593 3206
0 2 0 0 0 16 0 0 3 12 0 3
1329 2726
1329 3249
1496 3249
0 1 0 0 0 16 0 0 3 13 0 3
1299 2514
1299 3231
1496 3231
0 2 0 0 0 16 0 0 4 10 0 3
1261 2916
1261 3203
1495 3203
3 1 0 0 0 16 0 5 4 0 0 4
1403 3177
1467 3177
1467 3185
1495 3185
0 2 0 0 0 16 0 0 5 12 0 3
1152 2726
1152 3186
1354 3186
0 1 0 0 0 16 0 0 5 13 0 3
1202 2514
1202 3168
1354 3168
3 1 0 0 0 16 0 6 40 0 0 5
1665 2729
1690 2729
1690 175
1056 175
1056 80
3 2 0 0 0 16 0 9 6 0 0 4
946 2916
1603 2916
1603 2738
1616 2738
3 1 0 0 0 16 0 7 6 0 0 5
1644 2602
1644 2676
1600 2676
1600 2720
1616 2720
3 2 0 0 0 16 0 11 7 0 0 4
1090 2726
1567 2726
1567 2611
1595 2611
4 1 0 0 0 16 0 15 7 0 0 4
1153 2514
1566 2514
1566 2593
1595 2593
3 2 0 0 0 16 0 17 9 0 0 6
1396 2207
1511 2207
1511 3016
865 3016
865 2925
901 2925
1 0 0 0 0 16 0 8 0 0 88 8
758 2905
713 2905
713 2817
1546 2817
1546 419
477 419
477 405
461 405
2 1 0 0 0 16 0 8 9 0 0 3
794 2905
794 2907
901 2907
0 2 0 0 0 16 0 0 12 87 0 6
628 431
1478 431
1478 2846
881 2846
881 2770
927 2770
0 1 0 0 0 16 0 0 12 20 0 3
673 2669
673 2752
927 2752
0 2 0 0 0 16 0 0 13 91 0 4
557 436
28 436
28 2695
926 2695
1 0 0 0 0 16 0 10 0 0 29 4
711 2669
155 2669
155 195
303 195
2 1 0 0 0 16 0 10 13 0 0 4
747 2669
909 2669
909 2677
926 2677
3 2 0 0 0 16 0 12 11 0 0 4
972 2761
1013 2761
1013 2735
1044 2735
3 1 0 0 0 16 0 13 11 0 0 4
971 2686
1012 2686
1012 2717
1044 2717
2 3 0 0 0 16 0 14 15 0 0 4
933 2543
1098 2543
1098 2523
1108 2523
1 0 0 0 0 16 0 14 0 0 87 4
897 2543
19 2543
19 452
628 452
0 2 0 0 0 16 0 0 15 88 0 4
461 417
41 417
41 2514
1108 2514
3 1 0 0 0 16 0 16 15 0 0 4
1084 2434
1098 2434
1098 2505
1108 2505
2 0 0 0 0 16 0 16 0 0 91 4
1035 2443
58 2443
58 467
557 467
1 1 0 0 0 16 0 58 16 0 0 6
278 185
303 185
303 201
88 201
88 2425
1035 2425
3 2 0 0 0 16 0 18 17 0 0 4
1269 2245
1325 2245
1325 2216
1350 2216
3 1 0 0 0 16 0 19 17 0 0 4
1267 2175
1325 2175
1325 2198
1350 2198
0 2 0 0 0 16 0 0 18 36 0 4
1128 1806
734 1806
734 2254
1224 2254
0 1 0 0 0 16 0 0 18 42 0 5
1077 1600
1077 1641
840 1641
840 2236
1224 2236
0 2 0 0 0 16 0 0 19 39 0 3
1142 1928
1142 2184
1222 2184
3 1 0 0 0 16 0 20 19 0 0 4
1139 2152
1211 2152
1211 2166
1222 2166
0 2 0 0 0 16 0 0 20 41 0 5
1128 1730
1128 1847
815 1847
815 2161
1090 2161
0 1 0 0 0 16 0 0 20 42 0 5
1054 1600
1054 1654
1032 1654
1032 2143
1090 2143
3 1 0 0 0 16 0 21 41 0 0 5
1281 1944
1319 1944
1319 112
1094 112
1094 80
3 2 0 0 0 16 0 24 21 0 0 4
1032 1928
1154 1928
1154 1953
1232 1953
3 1 0 0 0 16 0 22 21 0 0 6
1234 1818
1254 1818
1254 1904
1193 1904
1193 1935
1232 1935
3 2 0 0 0 16 0 25 22 0 0 4
1121 1730
1151 1730
1151 1827
1185 1827
3 1 0 0 0 16 0 29 22 0 0 4
1029 1600
1168 1600
1168 1809
1185 1809
3 2 0 0 0 16 0 33 24 0 0 6
1109 1097
1140 1097
1140 1881
932 1881
932 1937
987 1937
2 1 0 0 0 16 0 23 24 0 0 4
901 1925
966 1925
966 1919
987 1919
0 1 0 0 0 16 0 0 23 88 0 4
461 429
114 429
114 1925
865 1925
3 2 0 0 0 16 0 27 25 0 0 4
1012 1776
1051 1776
1051 1739
1075 1739
3 1 0 0 0 16 0 28 25 0 0 4
1010 1697
1051 1697
1051 1721
1075 1721
0 2 0 0 0 16 0 0 27 87 0 4
628 472
135 472
135 1785
967 1785
0 1 0 0 0 16 0 0 27 59 0 4
431 230
158 230
158 1767
967 1767
0 2 0 0 0 16 0 0 28 91 0 4
557 477
170 477
170 1706
965 1706
2 1 0 0 0 16 0 26 28 0 0 4
802 1679
940 1679
940 1688
965 1688
0 1 0 0 0 16 0 0 26 59 0 4
431 210
196 210
196 1679
766 1679
1 2 0 0 0 16 0 63 29 0 0 8
392 79
433 79
433 150
352 150
352 263
216 263
216 1609
983 1609
4 1 0 0 0 16 0 31 29 0 0 4
908 1442
945 1442
945 1591
983 1591
2 3 0 0 0 16 0 30 31 0 0 4
670 1487
832 1487
832 1451
863 1451
0 1 0 0 0 16 0 0 30 87 0 4
628 484
232 484
232 1487
634 1487
0 2 0 0 0 16 0 0 31 88 0 4
461 459
244 459
244 1442
863 1442
3 1 0 0 0 16 0 32 31 0 0 4
782 1376
831 1376
831 1433
863 1433
1 2 0 0 0 16 0 59 32 0 0 6
387 187
431 187
431 310
279 310
279 1385
733 1385
0 1 0 0 0 16 0 0 32 91 0 4
557 494
309 494
309 1367
733 1367
3 2 0 0 0 16 0 34 33 0 0 4
1033 1134
1051 1134
1051 1106
1063 1106
3 1 0 0 0 16 0 35 33 0 0 4
1028 1066
1050 1066
1050 1088
1063 1088
0 2 0 0 0 16 0 0 34 72 0 6
970 684
983 684
983 781
698 781
698 1143
988 1143
0 1 0 0 0 16 0 0 34 73 0 4
969 629
826 629
826 1125
988 1125
0 2 0 0 0 16 0 0 35 70 0 7
982 837
982 884
1030 884
1030 1026
902 1026
902 1075
983 1075
3 1 0 0 0 16 0 36 35 0 0 6
986 976
1003 976
1003 1017
940 1017
940 1057
983 1057
0 2 0 0 0 16 0 0 36 72 0 5
959 699
959 913
871 913
871 985
937 985
0 1 0 0 0 16 0 0 36 73 0 6
969 610
946 610
946 925
897 925
897 967
937 967
3 1 0 0 0 16 0 37 42 0 0 5
1073 752
1158 752
1158 98
1134 98
1134 80
3 2 0 0 0 16 0 44 37 0 0 4
934 837
989 837
989 761
1024 761
3 1 0 0 0 16 0 38 37 0 0 6
1037 647
1048 647
1048 711
990 711
990 743
1024 743
3 2 0 0 0 16 0 45 38 0 0 4
942 699
970 699
970 656
988 656
3 1 0 0 0 16 0 49 38 0 0 4
944 593
969 593
969 638
988 638
2 2 0 0 0 16 0 43 44 0 0 4
815 852
877 852
877 846
889 846
0 1 0 0 0 16 0 0 43 88 0 4
461 442
410 442
410 852
779 852
1 1 0 0 0 16 0 53 44 0 0 4
718 389
752 389
752 828
889 828
3 2 0 0 0 16 0 47 45 0 0 4
740 744
872 744
872 708
896 708
3 1 0 0 0 16 0 48 45 0 0 4
744 655
872 655
872 690
896 690
0 2 0 0 0 16 0 0 47 87 0 4
628 502
473 502
473 753
695 753
0 1 0 0 0 16 0 0 47 90 0 4
525 319
333 319
333 735
695 735
0 2 0 0 0 16 0 0 48 91 0 4
557 512
510 512
510 664
699 664
2 1 0 0 0 16 0 46 48 0 0 4
591 649
683 649
683 646
699 646
0 1 0 0 0 16 0 0 46 90 0 4
525 328
353 328
353 649
555 649
1 2 0 0 0 16 0 64 49 0 0 4
494 77
852 77
852 602
898 602
4 1 0 0 0 16 0 51 49 0 0 4
844 579
872 579
872 584
898 584
2 3 0 0 0 16 0 50 51 0 0 4
639 603
771 603
771 588
799 588
1 1 0 0 0 16 0 56 50 0 0 6
614 403
628 403
628 562
581 562
581 603
603 603
1 2 0 0 0 16 0 54 51 0 0 4
435 399
461 399
461 579
799 579
3 1 0 0 0 16 0 52 51 0 0 4
725 530
770 530
770 570
799 570
1 2 0 0 0 16 0 60 52 0 0 6
498 185
525 185
525 340
385 340
385 539
676 539
1 1 0 0 0 16 0 55 52 0 0 4
535 402
557 402
557 521
676 521
19
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1596 3200 1633 3224
1606 3208 1622 3224
2 C2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1622 2711 1659 2735
1632 2719 1648 2735
2 F2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
905 2901 942 2925
915 2909 931 2925
2 Z2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1045 2708 1082 2732
1055 2716 1071 2732
2 Y2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1112 2497 1149 2521
1122 2505 1138 2521
2 X2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1352 2193 1389 2217
1362 2201 1378 2217
2 C1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1235 1927 1272 1951
1245 1935 1261 1951
2 F1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
990 1914 1027 1938
1000 1922 1016 1938
2 Z1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1078 1713 1115 1737
1088 1721 1104 1737
2 Y1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
986 1584 1023 1608
996 1592 1012 1608
2 X1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1066 1081 1103 1105
1076 1089 1092 1105
2 C0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1028 734 1065 758
1038 742 1054 758
2 F0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
995 13 1032 37
1005 21 1021 37
2 F3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1037 12 1074 36
1047 20 1063 36
2 F2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1073 14 1110 38
1083 22 1099 38
2 F1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1113 11 1150 35
1123 19 1139 35
2 F0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
893 823 930 847
903 831 919 847
2 Z0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
896 681 933 705
906 689 922 705
2 Y0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
899 577 936 601
909 585 925 601
2 X0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
