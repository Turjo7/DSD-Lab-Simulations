CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
50 900 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
42991634 0
0
6 Title:
5 Name:
0
0
0
59
13 Logic Switch~
5 610 736 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 Clear
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43564.7 0
0
13 Logic Switch~
5 609 774 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 CP
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
43564.7 1
0
13 Logic Switch~
5 124 961 0 10 11
0 46 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 I8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
43564.7 2
0
13 Logic Switch~
5 171 962 0 10 11
0 45 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 I7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
43564.7 3
0
13 Logic Switch~
5 266 963 0 1 11
0 43
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 I5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
43564.7 4
0
13 Logic Switch~
5 219 962 0 10 11
0 44 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 I6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
43564.7 5
0
14 Ascii Display~
172 3450 16 0 42 44
0 47 48 49 50 51 52 53 54 0
0 8224 8224 8224 8224 8224 8224 8224 8224 8224
8224 8224 8224 8224 8224 8224 8224 8224 8224 8224
8224 8224 8224 8224 8224 8224 8224 8224 8224 8224
8224 8224 8224
0
0 0 21088 0
4 1MEG
-15 -42 13 -34
5 DISP1
-3 -48 32 -40
0
0
102 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
%DE %5 0 %V
%DF %6 0 %V
%DG %7 0 %V
%DH %8 0 %V
0
0
0
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
82 0 0 512 1 0 0 0
4 DISP
8901 0 0
2
43564.7 6
0
5 4081~
219 1329 1493 0 3 22
0 4 3 2
0
0 0 624 0
4 4081
-7 -24 21 -16
5 T4out
-19 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 12 0
1 U
7361 0 0
2
43564.7 7
0
5 4081~
219 1338 1448 0 3 22
0 7 6 5
0
0 0 624 0
4 4081
-7 -24 21 -16
5 T6sub
-19 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 11 0
1 U
4747 0 0
2
43564.7 8
0
5 4081~
219 1339 1395 0 3 22
0 7 9 8
0
0 0 624 0
4 4081
-7 -24 21 -16
6 T6adSB
-22 -25 20 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 11 0
1 U
972 0 0
2
43564.7 9
0
5 4081~
219 1337 1345 0 3 22
0 11 9 10
0
0 0 624 0
4 4081
-7 -24 21 -16
6 T5adSB
-22 -25 20 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 11 0
1 U
3472 0 0
2
43564.7 10
0
5 4081~
219 1337 1303 0 3 22
0 4 3 12
0
0 0 624 0
4 4081
-7 -24 21 -16
5 T4dot
-19 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 11 0
1 U
9998 0 0
2
43564.7 11
0
5 4071~
219 1328 1252 0 3 22
0 16 15 14
0
0 0 624 0
4 4071
-7 -24 21 -16
4 T5T6
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 10 0
1 U
3536 0 0
2
43564.7 12
0
5 4081~
219 934 1274 0 3 22
0 7 9 15
0
0 0 624 0
4 4081
-7 -24 21 -16
6 T6adSB
-22 -25 20 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 9 0
1 U
4597 0 0
2
43564.7 13
0
5 4081~
219 931 1231 0 3 22
0 11 17 16
0
0 0 624 0
4 4081
-7 -24 21 -16
5 T5LDA
-19 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 9 0
1 U
3835 0 0
2
43564.7 14
0
5 4071~
219 1332 1112 0 3 22
0 19 20 13
0
0 0 624 0
4 4071
-7 -24 21 -16
4 T3T5
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 8 0
1 U
3670 0 0
2
43564.7 15
0
5 4081~
219 1008 1121 0 3 22
0 11 21 20
0
0 0 624 0
4 4081
-7 -24 21 -16
5 T5dot
-19 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 9 0
1 U
5616 0 0
2
43564.7 16
0
5 4071~
219 1336 1062 0 3 22
0 24 18 23
0
0 0 624 0
4 4071
-7 -24 21 -16
4 T1T4
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 8 0
1 U
9323 0 0
2
43564.7 17
0
5 4081~
219 1002 985 0 3 22
0 4 21 18
0
0 0 624 0
4 4081
-7 -24 21 -16
5 T4dot
-19 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 9 0
1 U
317 0 0
2
43564.7 18
0
14 Logic Display~
6 1278 814 0 1 2
10 24
0
0 0 53856 90
6 100MEG
3 -16 45 -8
2 T1
-9 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
43564.7 19
0
14 Logic Display~
6 1169 815 0 1 2
10 22
0
0 0 53856 90
6 100MEG
3 -16 45 -8
2 T2
-9 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
43564.7 20
0
14 Logic Display~
6 1061 809 0 1 2
10 19
0
0 0 53856 90
6 100MEG
3 -16 45 -8
2 T3
-9 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
43564.7 21
0
14 Logic Display~
6 942 812 0 1 2
10 4
0
0 0 53856 90
6 100MEG
3 -16 45 -8
2 T4
-9 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
43564.7 22
0
14 Logic Display~
6 824 811 0 1 2
10 11
0
0 0 53856 90
6 100MEG
3 -16 45 -8
2 T5
-9 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
43564.7 23
0
14 Logic Display~
6 695 812 0 1 2
10 7
0
0 0 53856 90
6 100MEG
3 -16 45 -8
2 T6
-9 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
43564.7 24
0
5 4071~
219 836 1042 0 3 22
0 17 9 21
0
0 0 624 0
4 4071
-7 -24 21 -16
6 LDadSB
-13 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 8 0
1 U
7100 0 0
2
43564.7 25
0
5 4071~
219 740 1092 0 3 22
0 6 25 9
0
0 0 624 0
4 4071
-7 -24 21 -16
6 ADDSUB
-13 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 8 0
1 U
3820 0 0
2
43564.7 26
0
14 Logic Display~
6 1422 1248 0 1 2
10 14
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 La
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
43564.7 27
0
14 Logic Display~
6 1423 1299 0 1 2
10 12
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 Ea
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
43564.7 28
0
14 Logic Display~
6 1421 1341 0 1 2
10 10
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 Lb
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
43564.7 29
0
14 Logic Display~
6 1423 1391 0 1 2
10 8
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 Eu
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
43564.7 30
0
14 Logic Display~
6 1425 1444 0 1 2
10 5
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 Su
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
43564.7 31
0
14 Logic Display~
6 1426 1489 0 1 2
10 2
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 Lo
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
43564.7 32
0
14 Logic Display~
6 1418 1195 0 1 2
10 18
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 Ei
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
43564.7 33
0
14 Logic Display~
6 1417 1155 0 1 2
10 19
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 Li
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9265 0 0
2
43564.7 34
0
14 Logic Display~
6 1415 1108 0 1 2
10 13
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 CE
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9442 0 0
2
43564.7 35
0
14 Logic Display~
6 1413 1058 0 1 2
10 23
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 Lm
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
43564.7 36
0
14 Logic Display~
6 1415 1016 0 1 2
10 24
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 Ep
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
43564.7 37
0
14 Logic Display~
6 1414 965 0 1 2
10 22
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 Cp
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
43564.7 38
0
6 JK RN~
219 777 667 0 6 22
0 11 28 27 29 33 7
0
0 0 4720 512
6 74LS73
-22 -42 20 -34
3 JK6
-13 -42 8 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 1 5 0
1 U
8464 0 0
2
43564.7 39
0
6 JK RN~
219 905 667 0 6 22
0 4 28 26 29 27 11
0
0 0 4720 512
6 74LS73
-22 -42 20 -34
3 JK5
-13 -42 8 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 2 5 0
1 U
7168 0 0
2
43564.7 40
0
6 JK RN~
219 1021 667 0 6 22
0 19 28 30 29 26 4
0
0 0 4720 512
6 74LS73
-22 -42 20 -34
3 JK4
-13 -42 8 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 1 6 0
1 U
3171 0 0
2
43564.7 41
0
6 JK RN~
219 1132 667 0 6 22
0 22 28 31 29 30 19
0
0 0 4720 512
6 74LS73
-22 -42 20 -34
3 JK3
-13 -42 8 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 2 6 0
1 U
4139 0 0
2
43564.7 42
0
6 JK RN~
219 1236 667 0 6 22
0 24 28 32 29 31 22
0
0 0 4720 512
6 74LS73
-22 -42 20 -34
3 JK2
-13 -42 8 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 1 7 0
1 U
6435 0 0
2
43564.7 43
0
6 JK RN~
219 1332 662 0 6 22
0 33 28 7 29 24 32
0
0 0 4720 512
6 74LS73
-22 -42 20 -34
3 JK1
-13 -42 8 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 2 7 0
1 U
5283 0 0
2
43564.7 44
0
5 4082~
219 453 1034 0 5 22
0 37 39 34 36 17
0
0 0 624 0
4 4082
-7 -24 21 -16
3 LDA
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
6874 0 0
2
43564.7 45
0
5 4082~
219 458 1105 0 5 22
0 40 39 34 36 25
0
0 0 624 0
4 4082
-7 -24 21 -16
3 ADD
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 1 0
1 U
5305 0 0
2
43564.7 46
0
5 4082~
219 461 1185 0 5 22
0 37 34 38 36 6
0
0 0 624 0
4 4082
-7 -24 21 -16
3 SUB
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
34 0 0
2
43564.7 47
0
5 4082~
219 466 1255 0 5 22
0 42 41 38 37 3
0
0 0 624 0
4 4082
-7 -24 21 -16
3 OUT
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
969 0 0
2
43564.7 48
0
5 4082~
219 471 1337 0 5 22
0 40 38 41 42 35
0
0 0 624 0
4 4082
-7 -24 21 -16
3 HLT
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
8402 0 0
2
43564.7 49
0
5 4041~
219 123 1025 0 3 22
0 46 36 42
0
0 0 112 270
4 4041
-14 -60 14 -52
2 A1
-7 -70 7 -62
0
15 DVDD=14;DGND=7;
41 %D [%14bi %7bi %1i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 6 5 4
10 9 8 13 12 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
3751 0 0
2
43564.7 50
0
5 4041~
219 174 1016 0 3 22
0 45 34 41
0
0 0 112 270
4 4041
-14 -60 14 -52
2 A2
-7 -70 7 -62
0
15 DVDD=14;DGND=7;
41 %D [%14bi %7bi %1i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 6 5 4 3 2 1 6 5 4
10 9 8 13 12 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
4292 0 0
2
43564.7 51
0
5 4041~
219 219 1012 0 3 22
0 44 39 38
0
0 0 112 270
4 4041
-14 -60 14 -52
2 A3
-7 -70 7 -62
0
15 DVDD=14;DGND=7;
41 %D [%14bi %7bi %1i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 3 2 1 6 5 4
10 9 8 13 12 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
6118 0 0
2
43564.7 52
0
5 4041~
219 267 1005 0 3 22
0 43 37 40
0
0 0 112 270
4 4041
-14 -60 14 -52
2 A4
-7 -70 7 -62
0
15 DVDD=14;DGND=7;
41 %D [%14bi %7bi %1i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 13 12 11 3 2 1 6 5 4
10 9 8 13 12 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
34 0 0
2
43564.7 53
0
14 Logic Display~
6 517 966 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 LDA
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6357 0 0
2
43564.7 54
0
14 Logic Display~
6 557 962 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 ADD
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
319 0 0
2
43564.7 55
0
14 Logic Display~
6 597 962 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 SUB
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3976 0 0
2
43564.7 56
0
14 Logic Display~
6 636 958 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 OUT
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7634 0 0
2
43564.7 57
0
14 Logic Display~
6 679 958 0 1 2
10 35
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 HLT
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
523 0 0
2
43564.7 58
0
99
3 1 2 0 0 4224 0 8 33 0 0 2
1350 1493
1410 1493
0 2 3 0 0 8192 0 0 8 14 0 3
636 1310
636 1502
1305 1502
0 1 4 0 0 8192 0 0 8 15 0 3
967 1294
967 1484
1305 1484
3 1 5 0 0 4224 0 9 32 0 0 2
1359 1448
1409 1448
0 2 6 0 0 8320 0 0 9 74 0 3
597 1185
597 1457
1314 1457
1 0 7 0 0 4096 0 9 0 0 8 3
1314 1439
712 1439
712 1386
1 3 8 0 0 4224 0 31 10 0 0 2
1407 1395
1360 1395
0 1 7 0 0 8192 0 0 10 45 0 3
712 1265
712 1386
1315 1386
0 2 9 0 0 8320 0 0 10 11 0 3
810 1352
810 1404
1315 1404
3 1 10 0 0 4224 0 11 30 0 0 2
1358 1345
1405 1345
0 2 9 0 0 0 0 0 11 20 0 3
810 1283
810 1354
1313 1354
0 1 11 0 0 8320 0 0 11 22 0 3
886 1222
886 1336
1313 1336
1 3 12 0 0 4224 0 29 12 0 0 2
1407 1303
1358 1303
0 2 3 0 0 8320 0 0 12 73 0 3
636 1253
636 1312
1313 1312
0 1 4 0 0 8320 0 0 12 42 0 3
967 976
967 1294
1313 1294
1 3 13 0 0 4224 0 36 16 0 0 2
1399 1112
1365 1112
1 3 14 0 0 4224 0 28 13 0 0 2
1406 1252
1361 1252
3 2 15 0 0 4224 0 14 13 0 0 4
955 1274
1290 1274
1290 1261
1315 1261
3 1 16 0 0 4224 0 15 13 0 0 4
952 1231
1288 1231
1288 1243
1315 1243
0 2 9 0 0 0 0 0 14 38 0 3
810 1051
810 1283
910 1283
0 2 17 0 0 4096 0 0 15 37 0 3
801 1033
801 1240
907 1240
1 0 11 0 0 0 0 15 0 0 65 3
907 1222
886 1222
886 884
0 1 18 0 0 8320 0 0 34 28 0 3
1059 985
1059 1199
1402 1199
1 0 19 0 0 4096 0 35 0 0 43 3
1401 1159
1077 1159
1077 1103
3 2 20 0 0 4224 0 17 16 0 0 2
1029 1121
1319 1121
0 2 21 0 0 4224 0 0 17 30 0 3
927 1042
927 1130
984 1130
1 0 22 0 0 16512 0 39 0 0 56 5
1398 969
1222 969
1222 876
1184 876
1184 650
3 2 18 0 0 0 0 19 18 0 0 4
1023 985
1272 985
1272 1071
1323 1071
1 3 23 0 0 4224 0 37 18 0 0 2
1397 1062
1369 1062
3 2 21 0 0 0 0 26 19 0 0 4
869 1042
955 1042
955 994
978 994
1 0 24 0 0 0 0 20 0 0 44 2
1293 817
1293 817
1 0 22 0 0 0 0 21 0 0 27 2
1184 818
1184 818
1 0 19 0 0 0 0 22 0 0 43 2
1076 812
1076 812
1 0 4 0 0 0 0 23 0 0 42 2
957 815
957 815
1 0 11 0 0 0 0 24 0 0 65 2
839 814
839 814
1 0 7 0 0 0 0 25 0 0 45 2
710 815
711 815
0 1 17 0 0 8320 0 0 26 76 0 3
517 1034
517 1033
823 1033
3 2 9 0 0 0 0 27 26 0 0 4
773 1092
788 1092
788 1051
823 1051
1 0 6 0 0 0 0 27 0 0 74 2
727 1083
597 1083
2 0 25 0 0 4224 0 27 0 0 75 2
727 1101
557 1101
0 1 24 0 0 8192 0 0 38 44 0 4
1293 868
1339 868
1339 1020
1399 1020
1 0 4 0 0 0 0 19 0 0 47 5
978 976
957 976
957 665
958 665
958 650
1 0 19 0 0 8320 0 16 0 0 52 3
1319 1103
1076 1103
1076 650
0 1 24 0 0 12416 0 0 18 60 0 5
1292 669
1292 697
1293 697
1293 1053
1323 1053
1 0 7 0 0 8192 0 14 0 0 64 4
910 1265
711 1265
711 649
730 649
5 3 26 0 0 4224 0 42 41 0 0 2
989 668
927 668
6 1 4 0 0 0 0 42 41 0 0 2
995 650
927 650
5 3 27 0 0 4224 0 41 40 0 0 2
873 668
799 668
0 2 28 0 0 4096 0 0 41 69 0 5
934 774
934 702
943 702
943 659
934 659
0 4 29 0 0 4096 0 0 41 70 0 2
903 736
903 698
5 3 30 0 0 4224 0 43 42 0 0 2
1100 668
1043 668
6 1 19 0 0 0 0 43 42 0 0 2
1106 650
1043 650
0 2 28 0 0 0 0 0 42 69 0 5
1050 774
1050 702
1059 702
1059 659
1050 659
0 4 29 0 0 0 0 0 42 70 0 2
1019 736
1019 698
5 3 31 0 0 4224 0 44 43 0 0 2
1204 668
1154 668
6 1 22 0 0 0 0 44 43 0 0 2
1210 650
1154 650
0 2 28 0 0 0 0 0 43 69 0 5
1161 774
1161 702
1170 702
1170 659
1161 659
0 4 29 0 0 0 0 0 43 70 0 2
1130 736
1130 698
6 3 32 0 0 8320 0 45 44 0 0 5
1306 645
1306 661
1279 661
1279 668
1258 668
1 5 24 0 0 0 0 44 45 0 0 6
1258 650
1292 650
1292 669
1292 669
1292 663
1300 663
0 2 28 0 0 0 0 0 44 69 0 5
1265 774
1265 702
1274 702
1274 659
1265 659
0 4 29 0 0 0 0 0 44 70 0 2
1234 736
1234 698
5 1 33 0 0 12416 0 40 45 0 0 6
745 668
742 668
742 595
1384 595
1384 645
1354 645
3 6 7 0 0 12416 0 45 40 0 0 6
1354 663
1365 663
1365 601
730 601
730 650
751 650
0 1 11 0 0 0 0 0 17 66 0 5
839 650
839 884
940 884
940 1112
984 1112
1 6 11 0 0 0 0 40 41 0 0 2
799 650
879 650
0 2 28 0 0 0 0 0 40 69 0 5
806 774
806 702
815 702
815 659
806 659
0 4 29 0 0 0 0 0 40 70 0 2
775 736
775 698
2 1 28 0 0 20608 0 45 2 0 0 6
1361 654
1382 654
1382 714
1383 714
1383 774
621 774
1 4 29 0 0 4224 0 1 45 0 0 5
622 736
1239 736
1239 735
1330 735
1330 693
0 2 34 0 0 4096 0 0 48 89 0 3
357 1039
357 1181
437 1181
5 1 35 0 0 8320 0 50 59 0 0 3
492 1337
679 1337
679 976
1 5 3 0 0 0 0 58 49 0 0 3
636 976
636 1255
487 1255
5 1 6 0 0 0 0 48 57 0 0 3
482 1185
597 1185
597 980
1 5 25 0 0 0 0 56 47 0 0 3
557 980
557 1105
479 1105
5 1 17 0 0 0 0 46 55 0 0 3
474 1034
517 1034
517 984
0 4 36 0 0 4096 0 0 48 88 0 3
369 1048
369 1199
437 1199
0 1 37 0 0 4096 0 0 48 91 0 3
347 1021
347 1172
437 1172
3 0 38 0 0 4096 0 48 0 0 97 2
437 1190
223 1190
0 4 36 0 0 0 0 0 47 88 0 3
325 1048
325 1119
434 1119
3 0 34 0 0 0 0 47 0 0 89 3
434 1110
313 1110
313 1039
0 2 39 0 0 8192 0 0 47 90 0 3
301 1030
301 1101
434 1101
1 0 40 0 0 4096 0 47 0 0 96 2
434 1092
271 1092
0 4 37 0 0 4224 0 0 49 91 0 3
287 1021
287 1269
442 1269
3 0 38 0 0 4096 0 49 0 0 97 2
442 1260
223 1260
2 0 41 0 0 4096 0 49 0 0 98 2
442 1251
178 1251
1 0 42 0 0 4096 0 49 0 0 99 2
442 1242
127 1242
4 2 36 0 0 4224 0 46 51 0 0 3
429 1048
118 1048
118 1041
3 2 34 0 0 4224 0 46 52 0 0 3
429 1039
169 1039
169 1032
2 2 39 0 0 8320 0 53 46 0 0 3
214 1028
214 1030
429 1030
2 1 37 0 0 0 0 54 46 0 0 2
262 1021
429 1021
1 1 43 0 0 8320 0 5 54 0 0 3
266 975
267 975
267 990
1 1 44 0 0 4224 0 6 53 0 0 2
219 974
219 997
1 1 45 0 0 8320 0 4 52 0 0 3
171 974
174 974
174 1001
1 1 46 0 0 8320 0 3 51 0 0 3
124 973
123 973
123 1010
3 1 40 0 0 4224 0 54 50 0 0 3
271 1021
271 1324
447 1324
3 2 38 0 0 4224 0 53 50 0 0 3
223 1028
223 1333
447 1333
3 3 41 0 0 4224 0 52 50 0 0 3
178 1032
178 1342
447 1342
3 4 42 0 0 8320 0 51 50 0 0 3
127 1041
127 1351
447 1351
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
