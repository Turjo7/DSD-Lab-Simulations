CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
39
13 Logic Switch~
5 28 742 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 31 33 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 201 1620 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 146 1621 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89878e-315 0
0
13 Logic Switch~
5 95 1623 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.89878e-315 0
0
7 Ground~
168 349 311 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5572 0 0
2
5.89878e-315 0
0
7 Ground~
168 423 626 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
5.89878e-315 0
0
7 Ground~
168 462 1509 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7361 0 0
2
5.89878e-315 0
0
2 +V
167 29 1368 0 1 3
0 4
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4747 0 0
2
5.89878e-315 0
0
2 +V
167 26 190 0 1 3
0 5
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
5.89878e-315 0
0
5 4049~
219 41 858 0 2 22
0 3 6
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U12E
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 12 0
1 U
3472 0 0
2
5.89878e-315 0
0
5 4049~
219 57 87 0 2 22
0 8 7
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U12D
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 12 0
1 U
9998 0 0
2
5.89878e-315 0
0
5 4049~
219 206 1515 0 2 22
0 9 12
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U12C
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 12 0
1 U
3536 0 0
2
5.89878e-315 0
0
5 4049~
219 155 1515 0 2 22
0 10 13
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U12B
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 12 0
1 U
4597 0 0
2
5.89878e-315 0
0
5 4049~
219 103 1516 0 2 22
0 11 15
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U12A
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 12 0
1 U
3835 0 0
2
5.89878e-315 0
0
14 Logic Display~
6 1098 1001 0 1 2
10 16
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.89878e-315 0
0
14 Logic Display~
6 1060 186 0 1 2
10 17
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.89878e-315 0
0
5 4071~
219 927 1006 0 3 22
0 19 18 16
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 11 0
1 U
9323 0 0
2
5.89878e-315 0
0
5 4071~
219 902 196 0 3 22
0 21 20 17
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 11 0
1 U
317 0 0
2
5.89878e-315 0
0
8 4-In OR~
219 745 1124 0 5 22
0 25 24 23 22 18
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U10B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
3108 0 0
2
5.89878e-315 0
0
8 4-In OR~
219 728 850 0 5 22
0 29 28 27 26 19
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U10A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
4299 0 0
2
5.89878e-315 0
0
8 4-In OR~
219 658 275 0 5 22
0 33 32 31 30 20
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U9B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 9 0
1 U
9672 0 0
2
5.89878e-315 0
0
8 4-In OR~
219 658 108 0 5 22
0 37 36 35 34 21
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U9A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 9 0
1 U
7876 0 0
2
5.89878e-315 0
0
5 4082~
219 271 1396 0 5 22
0 4 11 10 9 22
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 8 0
1 U
6369 0 0
2
5.89878e-315 0
0
5 4082~
219 270 1303 0 5 22
0 2 11 10 12 23
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 8 0
1 U
9172 0 0
2
5.89878e-315 0
0
5 4082~
219 271 1216 0 5 22
0 38 11 13 9 24
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U7B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 2 7 0
1 U
7100 0 0
2
5.89878e-315 0
0
5 4082~
219 273 1137 0 5 22
0 39 11 13 12 25
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U7A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 7 0
1 U
3820 0 0
2
5.89878e-315 0
0
5 4082~
219 274 1047 0 5 22
0 40 15 14 9 26
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U6B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 2 6 0
1 U
7678 0 0
2
5.89878e-315 0
0
5 4082~
219 275 962 0 5 22
0 2 15 10 12 27
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U6A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
961 0 0
2
5.89878e-315 0
0
5 4082~
219 277 883 0 5 22
0 6 15 13 9 28
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
3178 0 0
2
5.89878e-315 0
0
5 4082~
219 275 763 0 5 22
0 3 15 13 12 29
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
3409 0 0
2
5.89878e-315 0
0
5 4082~
219 274 568 0 5 22
0 5 11 10 9 30
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
3951 0 0
2
5.89878e-315 0
0
5 4082~
219 275 488 0 5 22
0 2 11 10 12 31
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
8885 0 0
2
5.89878e-315 0
0
5 4082~
219 275 414 0 5 22
0 41 11 13 9 32
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 2 3 0
1 U
3780 0 0
2
5.89878e-315 0
0
5 4082~
219 274 344 0 5 22
0 42 11 13 12 33
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 3 0
1 U
9265 0 0
2
5.89878e-315 0
0
5 4082~
219 274 263 0 5 22
0 2 15 10 9 34
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
9442 0 0
2
5.89878e-315 0
0
5 4082~
219 274 185 0 5 22
0 3 15 10 12 35
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
9424 0 0
2
5.89878e-315 0
0
5 4082~
219 274 115 0 5 22
0 7 15 13 9 36
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 1 0
1 U
9968 0 0
2
5.89878e-315 0
0
5 4082~
219 273 39 0 5 22
0 8 15 13 12 37
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
9281 0 0
2
5.89878e-315 0
0
86
1 1 2 0 0 8192 0 6 36 0 0 5
349 305
349 230
246 230
246 250
250 250
0 1 2 0 0 4224 0 0 29 5 0 5
355 1259
355 920
244 920
244 949
251 949
0 1 3 0 0 4224 0 0 37 12 0 3
69 719
69 172
250 172
1 1 2 0 0 0 0 7 33 0 0 5
423 620
423 450
242 450
242 475
251 475
1 1 2 0 0 0 0 8 25 0 0 5
462 1503
462 1259
232 1259
232 1290
246 1290
1 1 4 0 0 4224 0 9 24 0 0 3
29 1377
247 1377
247 1383
1 1 5 0 0 4224 0 10 32 0 0 4
26 199
26 546
250 546
250 555
2 1 6 0 0 12416 0 11 30 0 0 5
44 876
97 876
97 848
253 848
253 870
0 1 3 0 0 0 0 0 11 12 0 4
55 719
55 833
44 833
44 840
2 1 7 0 0 12416 0 12 38 0 0 5
60 105
86 105
86 95
250 95
250 102
0 1 8 0 0 4096 0 0 12 13 0 4
56 33
56 62
60 62
60 69
1 1 3 0 0 0 0 1 31 0 0 5
40 742
40 719
247 719
247 750
251 750
1 1 8 0 0 12416 0 2 39 0 0 4
43 33
86 33
86 26
249 26
0 4 9 0 0 4096 0 0 24 56 0 3
180 1429
247 1429
247 1410
0 3 10 0 0 4096 0 0 24 54 0 4
125 1412
236 1412
236 1401
247 1401
0 2 11 0 0 4096 0 0 24 49 0 4
78 1396
229 1396
229 1392
247 1392
0 4 12 0 0 4096 0 0 25 59 0 3
209 1351
246 1351
246 1317
0 3 10 0 0 4096 0 0 25 54 0 4
125 1329
242 1329
242 1308
246 1308
0 2 11 0 0 4096 0 0 25 49 0 4
78 1309
238 1309
238 1299
246 1299
0 4 9 0 0 0 0 0 26 56 0 3
180 1244
247 1244
247 1230
0 3 13 0 0 4096 0 0 26 60 0 4
158 1228
237 1228
237 1221
247 1221
0 2 11 0 0 0 0 0 26 49 0 4
78 1216
233 1216
233 1212
247 1212
0 4 12 0 0 4096 0 0 27 59 0 3
209 1190
249 1190
249 1151
0 3 13 0 0 4096 0 0 27 60 0 4
158 1157
238 1157
238 1142
249 1142
0 2 11 0 0 0 0 0 27 49 0 4
78 1149
228 1149
228 1133
249 1133
0 4 9 0 0 0 0 0 28 56 0 4
180 1116
245 1116
245 1061
250 1061
0 3 14 0 0 4224 0 0 28 0 0 4
128 1060
240 1060
240 1052
250 1052
0 2 15 0 0 4096 0 0 28 61 0 4
106 1047
240 1047
240 1043
250 1043
0 4 12 0 0 8192 0 0 29 59 0 3
209 975
209 976
251 976
0 3 10 0 0 4096 0 0 29 54 0 2
125 967
251 967
0 2 15 0 0 4096 0 0 29 61 0 3
106 954
251 954
251 958
0 4 9 0 0 0 0 0 30 56 0 4
180 902
247 902
247 897
253 897
0 3 13 0 0 8192 0 0 30 60 0 3
158 887
158 888
253 888
0 2 15 0 0 0 0 0 30 61 0 4
106 871
241 871
241 879
253 879
0 4 12 0 0 0 0 0 31 59 0 4
209 780
245 780
245 777
251 777
0 3 13 0 0 0 0 0 31 60 0 4
158 759
223 759
223 768
251 768
0 2 15 0 0 0 0 0 31 61 0 4
106 743
231 743
231 759
251 759
0 4 9 0 0 0 0 0 32 56 0 4
180 600
237 600
237 582
250 582
0 3 10 0 0 0 0 0 32 54 0 4
125 576
236 576
236 573
250 573
0 2 11 0 0 4096 0 0 32 49 0 4
78 559
243 559
243 564
250 564
0 4 12 0 0 0 0 0 33 59 0 4
209 525
243 525
243 502
251 502
0 3 10 0 0 0 0 0 33 54 0 4
125 508
235 508
235 493
251 493
0 2 11 0 0 0 0 0 33 49 0 4
78 492
226 492
226 484
251 484
0 4 9 0 0 0 0 0 34 56 0 4
180 434
246 434
246 428
251 428
0 3 13 0 0 0 0 0 34 60 0 3
158 417
158 419
251 419
0 2 11 0 0 8192 0 0 34 49 0 3
78 411
78 410
251 410
0 4 12 0 0 0 0 0 35 59 0 3
209 362
250 362
250 358
0 3 13 0 0 0 0 0 35 60 0 4
158 350
239 350
239 349
250 349
0 2 11 0 0 8320 0 0 35 64 0 4
107 1564
78 1564
78 340
250 340
0 4 9 0 0 0 0 0 36 56 0 4
180 280
243 280
243 277
250 277
0 3 10 0 0 0 0 0 36 54 0 3
125 265
125 268
250 268
0 2 15 0 0 0 0 0 36 61 0 3
106 260
106 259
250 259
0 4 12 0 0 0 0 0 37 59 0 4
209 223
246 223
246 199
250 199
0 3 10 0 0 8320 0 0 37 63 0 6
166 1567
125 1567
125 203
237 203
237 190
250 190
0 2 15 0 0 0 0 0 37 61 0 4
106 192
231 192
231 181
250 181
0 4 9 0 0 8320 0 0 38 62 0 5
237 1548
180 1548
180 141
250 141
250 129
0 3 13 0 0 0 0 0 38 60 0 4
158 131
227 131
227 120
250 120
0 2 15 0 0 0 0 0 38 61 0 3
106 112
106 111
250 111
2 4 12 0 0 4224 0 13 39 0 0 3
209 1497
209 53
249 53
2 3 13 0 0 4224 0 14 39 0 0 3
158 1497
158 44
249 44
2 2 15 0 0 4224 0 15 39 0 0 3
106 1498
106 35
249 35
1 1 9 0 0 0 0 3 13 0 0 5
213 1620
237 1620
237 1538
209 1538
209 1533
1 1 10 0 0 0 0 4 14 0 0 5
158 1621
166 1621
166 1538
158 1538
158 1533
1 1 11 0 0 0 0 5 15 0 0 4
107 1623
107 1539
106 1539
106 1534
3 1 16 0 0 8320 0 18 16 0 0 3
960 1006
960 1005
1082 1005
3 1 17 0 0 4224 0 19 17 0 0 4
935 196
1026 196
1026 190
1044 190
5 2 18 0 0 8320 0 20 18 0 0 4
778 1124
886 1124
886 1015
914 1015
5 1 19 0 0 8320 0 21 18 0 0 4
761 850
886 850
886 997
914 997
5 2 20 0 0 4224 0 22 19 0 0 4
691 275
868 275
868 205
889 205
5 1 21 0 0 4224 0 23 19 0 0 4
691 108
868 108
868 187
889 187
5 4 22 0 0 4224 0 24 20 0 0 4
292 1396
702 1396
702 1138
728 1138
5 3 23 0 0 4224 0 25 20 0 0 4
291 1303
674 1303
674 1129
728 1129
5 2 24 0 0 4224 0 26 20 0 0 4
292 1216
652 1216
652 1120
728 1120
5 1 25 0 0 4224 0 27 20 0 0 4
294 1137
643 1137
643 1111
728 1111
5 4 26 0 0 4224 0 28 21 0 0 4
295 1047
658 1047
658 864
711 864
5 3 27 0 0 4224 0 29 21 0 0 4
296 962
637 962
637 855
711 855
5 2 28 0 0 4224 0 30 21 0 0 4
298 883
615 883
615 846
711 846
5 1 29 0 0 4224 0 31 21 0 0 4
296 763
689 763
689 837
711 837
5 4 30 0 0 4224 0 32 22 0 0 5
295 568
658 568
658 300
641 300
641 289
5 3 31 0 0 4224 0 33 22 0 0 4
296 488
636 488
636 280
641 280
5 2 32 0 0 4224 0 34 22 0 0 4
296 414
628 414
628 271
641 271
5 1 33 0 0 4224 0 35 22 0 0 4
295 344
619 344
619 262
641 262
5 4 34 0 0 4224 0 36 23 0 0 7
295 263
596 263
596 200
648 200
648 138
641 138
641 122
5 3 35 0 0 4224 0 37 23 0 0 6
295 185
632 185
632 119
637 119
637 113
641 113
5 2 36 0 0 4224 0 38 23 0 0 4
295 115
630 115
630 104
641 104
5 1 37 0 0 4224 0 39 23 0 0 4
294 39
629 39
629 95
641 95
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
