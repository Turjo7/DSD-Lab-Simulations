CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 326 288 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
7 Jswitch
-23 -26 26 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43548.4 0
0
13 Logic Switch~
5 646 515 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 P5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43548.4 0
0
13 Logic Switch~
5 142 313 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 P4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 0 0 -1 0
1 V
3124 0 0
2
43548.4 0
0
13 Logic Switch~
5 208 357 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
7 KSwitch
-23 -26 26 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43548.4 0
0
13 Logic Switch~
5 174 499 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
5 clock
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43548.4 0
0
14 Logic Display~
6 849 273 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
43548.4 0
0
7 Pulser~
4 500 508 0 11 12
0 5 9 7 10 0 0 5 5 -1
7 1
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
8901 0 0
2
43548.4 0
0
6 JK RN~
219 671 356 0 6 22
0 6 7 4 2 11 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
7361 0 0
2
43548.4 0
0
6
1 4 2 0 0 8320 0 2 8 0 0 3
658 515
671 515
671 387
6 1 3 0 0 4224 0 8 6 0 0 4
695 339
798 339
798 291
849 291
3 1 4 0 0 4224 0 8 4 0 0 2
647 357
220 357
1 1 5 0 0 4224 0 7 5 0 0 2
476 499
186 499
1 1 6 0 0 4224 0 8 1 0 0 4
647 339
389 339
389 288
338 288
3 2 7 0 0 8320 0 7 8 0 0 4
524 499
588 499
588 348
640 348
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
