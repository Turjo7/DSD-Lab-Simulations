CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 464 108 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43509.5 0
0
13 Logic Switch~
5 401 110 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43509.5 0
0
13 Logic Switch~
5 347 105 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43509.5 0
0
13 Logic Switch~
5 283 106 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43509.5 0
0
13 Logic Switch~
5 223 114 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 Bi
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43509.5 0
0
13 Logic Switch~
5 156 120 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 Ai
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
43509.5 0
0
5 4081~
219 948 468 0 3 22
0 4 3 2
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
8901 0 0
2
43509.5 0
0
14 Logic Display~
6 1063 336 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
43509.5 0
0
14 Logic Display~
6 998 208 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
43509.5 0
0
5 4071~
219 1035 462 0 3 22
0 7 2 5
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
972 0 0
2
43509.5 0
0
5 4030~
219 850 509 0 3 22
0 9 8 3
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
3472 0 0
2
43509.5 0
0
5 4081~
219 850 449 0 3 22
0 9 8 7
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
9998 0 0
2
43509.5 0
0
5 4070~
219 916 225 0 3 22
0 10 4 6
0
0 0 624 0
4 4070
-7 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
3536 0 0
2
43509.5 0
0
5 4070~
219 850 214 0 3 22
0 9 8 10
0
0 0 624 0
4 4070
-7 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
4597 0 0
2
43509.5 0
0
5 4081~
219 578 411 0 3 22
0 12 11 4
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
3835 0 0
2
43509.5 0
0
5 4049~
219 309 125 0 2 22
0 13 12
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
3670 0 0
2
43509.5 0
0
5 4049~
219 252 140 0 2 22
0 15 14
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
5616 0 0
2
43509.5 0
0
5 4071~
219 638 320 0 3 22
0 19 18 8
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
9323 0 0
2
43509.5 0
0
5 4081~
219 577 349 0 3 22
0 16 14 18
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
317 0 0
2
43509.5 0
0
5 4081~
219 575 299 0 3 22
0 15 17 19
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
3108 0 0
2
43509.5 0
0
5 4071~
219 702 206 0 3 22
0 21 20 9
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
4299 0 0
2
43509.5 0
0
5 4081~
219 637 204 0 3 22
0 23 22 21
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
9672 0 0
2
43509.5 0
0
5 4049~
219 427 124 0 2 22
0 17 24
0
0 0 624 270
4 4049
-7 -24 21 -16
3 U3A
16 -8 37 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
7876 0 0
2
43509.5 0
0
5 4081~
219 569 234 0 3 22
0 13 24 22
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
6369 0 0
2
43509.5 0
0
5 4030~
219 559 180 0 3 22
0 16 15 23
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
9172 0 0
2
43509.5 0
0
35
3 2 2 0 0 8320 0 7 10 0 0 3
969 468
969 471
1022 471
2 0 3 0 0 4096 0 7 0 0 8 2
924 477
923 477
1 0 4 0 0 0 0 7 0 0 7 2
924 459
924 459
3 1 5 0 0 4224 0 10 8 0 0 3
1068 462
1068 354
1063 354
3 1 6 0 0 8320 0 13 9 0 0 3
949 225
949 226
998 226
3 1 7 0 0 12416 0 12 10 0 0 6
871 449
893 449
893 435
989 435
989 453
1022 453
0 0 4 0 0 4096 0 0 0 13 0 3
897 411
897 459
930 459
3 0 3 0 0 4224 0 11 0 0 0 4
883 509
923 509
923 477
930 477
2 0 8 0 0 4096 0 11 0 0 11 3
834 518
701 518
701 458
1 0 9 0 0 4096 0 11 0 0 12 3
834 500
743 500
743 440
2 0 8 0 0 8320 0 12 0 0 15 3
826 458
701 458
701 320
1 0 9 0 0 8320 0 12 0 0 16 3
826 440
743 440
743 205
3 2 4 0 0 4224 0 15 13 0 0 3
599 411
900 411
900 234
1 3 10 0 0 8320 0 13 14 0 0 3
900 216
900 214
883 214
3 2 8 0 0 0 0 18 14 0 0 4
671 320
734 320
734 223
834 223
3 1 9 0 0 0 0 21 14 0 0 3
735 206
735 205
834 205
1 2 11 0 0 4224 0 1 15 0 0 3
476 108
476 420
554 420
2 1 12 0 0 4224 0 16 15 0 0 3
330 125
330 402
554 402
1 0 13 0 0 4096 0 16 0 0 33 2
294 125
295 125
2 2 14 0 0 8320 0 17 19 0 0 3
273 140
273 358
553 358
1 0 15 0 0 4096 0 17 0 0 34 2
237 140
235 140
0 1 16 0 0 8320 0 0 19 35 0 3
359 171
359 340
553 340
1 2 17 0 0 4224 0 2 20 0 0 3
413 110
413 308
551 308
0 1 15 0 0 8320 0 0 20 34 0 3
235 189
235 290
551 290
3 2 18 0 0 8320 0 19 18 0 0 4
598 349
610 349
610 329
625 329
3 1 19 0 0 4224 0 20 18 0 0 4
596 299
613 299
613 311
625 311
1 2 20 0 0 8320 0 6 21 0 0 5
168 120
168 258
680 258
680 215
689 215
3 1 21 0 0 4224 0 22 21 0 0 3
658 204
689 204
689 197
3 2 22 0 0 8320 0 24 22 0 0 4
590 234
606 234
606 213
613 213
3 1 23 0 0 8320 0 25 22 0 0 4
592 180
605 180
605 195
613 195
2 2 24 0 0 8320 0 23 24 0 0 3
430 142
430 243
545 243
1 1 17 0 0 0 0 2 23 0 0 3
413 110
413 106
430 106
1 1 13 0 0 8320 0 4 24 0 0 3
295 106
295 225
545 225
1 2 15 0 0 0 0 5 25 0 0 3
235 114
235 189
543 189
1 1 16 0 0 0 0 25 3 0 0 3
543 171
359 171
359 105
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
