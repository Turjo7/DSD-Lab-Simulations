CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1950 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
3 100 1 2 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
67
13 Logic Switch~
5 45 1127 0 1 11
0 38
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 I7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89888e-315 0
0
13 Logic Switch~
5 122 1129 0 1 11
0 37
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 I6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89888e-315 0
0
13 Logic Switch~
5 207 1131 0 1 11
0 36
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 I5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89888e-315 0
0
13 Logic Switch~
5 284 1133 0 1 11
0 35
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 I4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89888e-315 0
0
13 Logic Switch~
5 693 885 0 10 11
0 45 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 CP
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.89888e-315 5.26354e-315
0
13 Logic Switch~
5 694 847 0 10 11
0 46 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 Clear
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.89888e-315 0
0
5 4049~
219 960 2290 0 2 22
0 3 2
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 16 0
1 U
8901 0 0
2
5.89888e-315 0
0
5 4081~
219 891 2288 0 3 22
0 5 4 3
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U10B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 18 0
1 U
7361 0 0
2
5.89888e-315 0
0
5 4049~
219 992 2143 0 2 22
0 7 6
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 16 0
1 U
4747 0 0
2
5.89888e-315 0
0
5 4081~
219 914 2143 0 3 22
0 9 8 7
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 18 0
1 U
972 0 0
2
5.89888e-315 0
0
5 4081~
219 906 2030 0 3 22
0 9 11 10
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 17 0
1 U
3472 0 0
2
5.89888e-315 0
0
5 4081~
219 131 680 0 3 22
0 11 13 12
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 17 0
1 U
9998 0 0
2
5.89888e-315 0
0
5 4081~
219 652 637 0 3 22
0 5 4 14
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 17 0
1 U
3536 0 0
2
5.89888e-315 0
0
5 4049~
219 1098 1842 0 2 22
0 16 15
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 16 0
1 U
4597 0 0
2
5.89888e-315 0
0
5 4071~
219 1019 1848 0 3 22
0 18 17 16
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 15 0
1 U
3835 0 0
2
5.89888e-315 0
0
5 4081~
219 914 1908 0 3 22
0 9 11 17
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 17 0
1 U
3670 0 0
2
5.89888e-315 0
0
5 4071~
219 813 1880 0 3 22
0 19 13 9
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 15 0
1 U
5616 0 0
2
5.89888e-315 0
0
5 4081~
219 828 1784 0 3 22
0 8 20 18
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 14 0
1 U
9323 0 0
2
5.89888e-315 0
0
5 4049~
219 900 1694 0 2 22
0 22 21
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 16 0
1 U
317 0 0
2
5.89888e-315 0
0
5 4081~
219 829 1694 0 3 22
0 23 5 22
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 14 0
1 U
3108 0 0
2
5.89888e-315 0
0
5 4049~
219 475 612 0 2 22
0 25 24
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 16 0
1 U
4299 0 0
2
5.89888e-315 0
0
5 4049~
219 1016 1557 0 2 22
0 27 26
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U1F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 9 0
1 U
9672 0 0
2
5.89888e-315 0
0
5 4071~
219 941 1558 0 3 22
0 28 25 27
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 15 0
1 U
7876 0 0
2
5.89888e-315 0
0
5 4081~
219 877 1519 0 3 22
0 23 8 28
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 14 0
1 U
6369 0 0
2
5.89888e-315 0
0
5 4049~
219 1051 1445 0 2 22
0 30 29
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U1E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 9 0
1 U
9172 0 0
2
5.89888e-315 0
0
5 4071~
219 974 1446 0 3 22
0 32 31 30
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 15 0
1 U
7100 0 0
2
5.89888e-315 0
0
5 4081~
219 918 1418 0 3 22
0 23 5 32
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 14 0
1 U
3820 0 0
2
5.89888e-315 0
0
8 3-In OR~
219 815 1397 0 4 22
0 20 19 13 23
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 13 0
1 U
7678 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 845 437 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L23
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 800 440 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L22
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 747 441 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L21
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 692 442 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L20
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 527 443 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L19
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 474 443 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L18
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 423 442 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L17
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9265 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 371 444 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L16
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9442 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 240 448 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 186 449 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 137 450 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 87 451 0 1 2
10 33
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 386 1066 0 1 2
10 34
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 453 1068 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 514 1069 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 578 1069 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6435 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 630 1069 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
5.89888e-315 0
0
5 4082~
219 440 1795 0 5 22
0 35 36 37 38 34
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 12 0
1 U
6874 0 0
2
5.89888e-315 0
0
5 4082~
219 440 1674 0 5 22
0 39 36 37 38 4
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 11 0
1 U
5305 0 0
2
5.89888e-315 0
0
5 4082~
219 441 1550 0 5 22
0 39 36 41 40 13
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 11 0
1 U
34 0 0
2
5.89888e-315 0
0
5 4082~
219 441 1424 0 5 22
0 35 42 41 40 19
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
969 0 0
2
5.89888e-315 0
0
5 4082~
219 443 1298 0 5 22
0 39 42 41 40 20
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
8402 0 0
2
5.89888e-315 0
0
5 4049~
219 52 1216 0 2 22
0 38 40
0
0 0 624 270
4 4049
-7 -24 21 -16
3 U1D
16 -8 37 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 9 0
1 U
3751 0 0
2
5.89888e-315 0
0
5 4049~
219 137 1212 0 2 22
0 37 41
0
0 0 624 270
4 4049
-7 -24 21 -16
3 U1C
16 -8 37 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 9 0
1 U
4292 0 0
2
5.89888e-315 0
0
5 4049~
219 217 1206 0 2 22
0 36 42
0
0 0 624 270
4 4049
-7 -24 21 -16
3 U1B
16 -8 37 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 9 0
1 U
6118 0 0
2
5.89888e-315 0
0
5 4049~
219 293 1207 0 2 22
0 35 39
0
0 0 624 270
4 4049
-7 -24 21 -16
3 U1A
16 -8 37 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 9 0
1 U
34 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 532 720 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6357 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 218 731 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
319 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 285 729 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3976 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 337 728 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7634 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 411 727 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
523 0 0
2
5.89888e-315 0
0
14 Logic Display~
6 475 727 0 1 2
10 33
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
5.89888e-315 0
0
6 JK RN~
219 1416 773 0 6 22
0 50 45 11 46 31 49
0
0 0 4720 512
6 74LS73
-22 -42 20 -34
4 JK3B
-16 -42 12 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 2 8 0
1 U
6901 0 0
2
5.89888e-315 5.32571e-315
0
6 JK RN~
219 1320 778 0 6 22
0 31 45 49 46 48 33
0
0 0 4720 512
6 74LS73
-22 -42 20 -34
4 JK3A
-16 -42 12 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 1 8 0
1 U
842 0 0
2
5.89888e-315 5.30499e-315
0
6 JK RN~
219 1216 778 0 6 22
0 33 45 48 46 47 25
0
0 0 4720 512
6 74LS73
-22 -42 20 -34
4 JK2B
-16 -42 12 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 2 7 0
1 U
3277 0 0
2
5.89888e-315 5.26354e-315
0
6 JK RN~
219 1105 778 0 6 22
0 25 45 47 46 43 5
0
0 0 4720 512
6 74LS73
-22 -42 20 -34
4 JK2A
-16 -42 12 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 1 7 0
1 U
4212 0 0
2
5.89888e-315 0
0
6 JK RN~
219 989 778 0 6 22
0 5 45 43 46 44 8
0
0 0 4720 512
6 74LS73
-22 -42 20 -34
4 JK1B
-16 -42 12 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 2 6 0
1 U
4720 0 0
2
5.89888e-315 5.48113e-315
0
6 JK RN~
219 861 778 0 6 22
0 8 45 44 46 50 11
0
0 0 4720 512
6 74LS73
-22 -42 20 -34
4 JK1A
-16 -42 12 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 1 6 0
1 U
5551 0 0
2
5.89888e-315 5.47984e-315
0
14 Ascii Display~
172 3534 127 0 42 44
0 51 52 53 54 55 56 57 58 0
0 8224 8224 8224 8224 8224 8224 8224 8224 8224
8224 8224 8224 8224 8224 8224 8224 8224 8224 8224
8224 8224 8224 8224 8224 8224 8224 8224 8224 8224
8224 8224 8224
0
0 0 21088 0
4 1MEG
-15 -42 13 -34
5 DISP1
-3 -48 32 -40
0
0
102 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
%DE %5 0 %V
%DF %6 0 %V
%DG %7 0 %V
%DH %8 0 %V
0
0
0
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
82 0 0 512 1 0 0 0
4 DISP
6986 0 0
2
5.89888e-315 5.36716e-315
0
109
2 1 2 0 0 8320 0 7 29 0 0 5
981 2290
1819 2290
1819 465
845 465
845 455
3 1 3 0 0 8320 0 8 7 0 0 3
912 2288
912 2290
945 2290
0 2 4 0 0 8320 0 0 8 52 0 4
508 1138
495 1138
495 2297
867 2297
0 1 5 0 0 8320 0 0 8 82 0 4
337 782
315 782
315 2279
867 2279
2 1 6 0 0 8320 0 9 30 0 0 5
1013 2143
1767 2143
1767 476
800 476
800 458
3 1 7 0 0 4224 0 10 9 0 0 2
935 2143
977 2143
0 2 8 0 0 16512 0 0 10 81 0 6
285 884
258 884
258 913
848 913
848 2152
890 2152
0 1 9 0 0 4096 0 0 10 11 0 3
867 2021
867 2134
890 2134
3 1 10 0 0 8320 0 11 31 0 0 5
927 2030
1711 2030
1711 501
747 501
747 459
0 2 11 0 0 12288 0 0 11 14 0 5
218 804
218 984
736 984
736 2039
882 2039
0 1 9 0 0 4224 0 0 11 23 0 3
852 1880
852 2021
882 2021
3 1 12 0 0 12416 0 12 32 0 0 5
152 680
175 680
175 481
692 481
692 460
0 2 13 0 0 24576 0 0 12 53 0 10
528 1157
417 1157
417 1137
345 1137
345 1077
105 1077
105 708
79 708
79 689
107 689
0 1 11 0 0 0 0 0 12 80 0 5
245 752
245 804
42 804
42 671
107 671
3 1 14 0 0 8320 0 13 33 0 0 7
673 637
685 637
685 496
575 496
575 466
527 466
527 461
0 2 4 0 0 0 0 0 13 52 0 6
508 1186
568 1186
568 1098
553 1098
553 646
628 646
0 1 5 0 0 0 0 0 13 82 0 4
337 807
607 807
607 628
628 628
2 1 15 0 0 8320 0 14 34 0 0 7
1119 1842
1681 1842
1681 515
561 515
561 489
474 489
474 461
3 1 16 0 0 4224 0 15 14 0 0 4
1052 1848
1072 1848
1072 1842
1083 1842
3 2 17 0 0 8320 0 16 15 0 0 4
935 1908
985 1908
985 1857
1006 1857
3 1 18 0 0 4224 0 18 15 0 0 4
849 1784
968 1784
968 1839
1006 1839
0 2 11 0 0 4224 0 0 16 80 0 3
649 752
649 1917
890 1917
3 1 9 0 0 0 0 17 16 0 0 4
846 1880
876 1880
876 1899
890 1899
0 2 13 0 0 8320 0 0 17 53 0 4
528 1138
548 1138
548 1889
800 1889
0 1 19 0 0 8320 0 0 17 54 0 4
578 1123
598 1123
598 1871
800 1871
0 2 20 0 0 4224 0 0 18 48 0 3
645 1101
645 1793
804 1793
0 1 8 0 0 0 0 0 18 81 0 3
663 993
663 1775
804 1775
2 1 21 0 0 12416 0 19 35 0 0 5
921 1694
1637 1694
1637 528
423 528
423 460
3 1 22 0 0 4224 0 20 19 0 0 2
850 1694
885 1694
0 2 5 0 0 0 0 0 20 82 0 3
679 969
679 1703
805 1703
0 1 23 0 0 8320 0 0 20 39 0 4
855 1442
779 1442
779 1685
805 1685
2 1 24 0 0 12416 0 21 36 0 0 5
496 612
540 612
540 506
371 506
371 462
0 1 25 0 0 8192 0 0 21 83 0 4
411 785
444 785
444 612
460 612
2 1 26 0 0 12416 0 22 37 0 0 5
1037 1557
1608 1557
1608 542
240 542
240 466
3 1 27 0 0 8320 0 23 22 0 0 3
974 1558
974 1557
1001 1557
0 2 25 0 0 4096 0 0 23 83 0 3
706 956
706 1567
928 1567
3 1 28 0 0 8320 0 24 23 0 0 4
898 1519
908 1519
908 1549
928 1549
0 2 8 0 0 0 0 0 24 81 0 3
758 993
758 1528
853 1528
0 1 23 0 0 0 0 0 24 45 0 5
855 1397
855 1489
820 1489
820 1510
853 1510
2 1 29 0 0 12416 0 25 38 0 0 5
1072 1445
1589 1445
1589 557
186 557
186 467
3 1 30 0 0 8320 0 26 25 0 0 3
1007 1446
1007 1445
1036 1445
0 2 31 0 0 4096 0 0 26 85 0 5
808 925
808 1364
717 1364
717 1455
961 1455
3 1 32 0 0 8320 0 27 26 0 0 4
939 1418
954 1418
954 1437
961 1437
0 2 5 0 0 0 0 0 27 82 0 3
786 969
786 1427
894 1427
4 1 23 0 0 0 0 28 27 0 0 4
848 1397
887 1397
887 1409
894 1409
0 3 13 0 0 0 0 0 28 53 0 6
528 1117
560 1117
560 1191
692 1191
692 1406
802 1406
0 2 19 0 0 0 0 0 28 54 0 4
578 1108
605 1108
605 1397
803 1397
0 1 20 0 0 0 0 0 28 55 0 4
630 1101
751 1101
751 1388
802 1388
0 1 31 0 0 24704 0 0 39 85 0 8
826 925
826 1232
1038 1232
1038 1229
1564 1229
1564 569
137 569
137 468
0 1 33 0 0 24704 0 0 40 84 0 8
876 944
876 1161
1038 1161
1038 1153
1548 1153
1548 580
87 580
87 469
1 5 34 0 0 12416 0 41 46 0 0 5
386 1084
386 1119
483 1119
483 1795
461 1795
5 1 4 0 0 0 0 47 42 0 0 7
461 1674
508 1674
508 1111
489 1111
489 1095
453 1095
453 1086
5 1 13 0 0 0 0 48 43 0 0 5
462 1550
528 1550
528 1098
514 1098
514 1087
5 1 19 0 0 0 0 49 44 0 0 3
462 1424
578 1424
578 1087
5 1 20 0 0 0 0 50 45 0 0 3
464 1298
630 1298
630 1087
0 1 35 0 0 8320 0 0 46 71 0 4
387 1229
367 1229
367 1782
416 1782
0 2 36 0 0 8192 0 0 46 62 0 3
277 1670
277 1791
416 1791
0 3 37 0 0 8192 0 0 46 61 0 3
209 1679
209 1800
416 1800
0 4 38 0 0 8192 0 0 46 60 0 3
149 1688
149 1809
416 1809
0 4 38 0 0 8320 0 0 47 76 0 4
77 1177
7 1177
7 1688
416 1688
0 3 37 0 0 8320 0 0 47 77 0 4
159 1169
187 1169
187 1679
416 1679
0 2 36 0 0 8320 0 0 47 66 0 4
272 1260
252 1260
252 1670
416 1670
0 1 39 0 0 4224 0 0 47 75 0 3
347 1285
347 1661
416 1661
0 4 40 0 0 12416 0 0 48 72 0 4
55 1267
20 1267
20 1564
417 1564
0 3 41 0 0 12416 0 0 48 73 0 4
140 1257
84 1257
84 1555
417 1555
0 2 36 0 0 0 0 0 48 78 0 4
232 1168
272 1168
272 1546
417 1546
0 1 39 0 0 0 0 0 48 75 0 3
322 1285
322 1537
417 1537
0 4 40 0 0 0 0 0 49 72 0 4
55 1282
35 1282
35 1438
417 1438
0 3 41 0 0 0 0 0 49 73 0 4
140 1283
110 1283
110 1429
417 1429
0 2 42 0 0 12416 0 0 49 74 0 4
220 1279
204 1279
204 1420
417 1420
0 1 35 0 0 0 0 0 49 79 0 4
323 1164
387 1164
387 1411
417 1411
2 4 40 0 0 0 0 51 50 0 0 3
55 1234
55 1312
419 1312
2 3 41 0 0 0 0 52 50 0 0 3
140 1230
140 1303
419 1303
2 2 42 0 0 0 0 53 50 0 0 5
220 1224
220 1296
356 1296
356 1294
419 1294
2 1 39 0 0 0 0 54 50 0 0 3
296 1225
296 1285
419 1285
1 1 38 0 0 0 0 1 51 0 0 5
57 1127
77 1127
77 1190
55 1190
55 1198
1 1 37 0 0 0 0 2 52 0 0 5
134 1129
159 1129
159 1180
140 1180
140 1194
1 1 36 0 0 0 0 3 53 0 0 5
219 1131
232 1131
232 1173
220 1173
220 1188
1 1 35 0 0 0 0 4 54 0 0 5
296 1133
323 1133
323 1171
296 1171
296 1189
0 1 11 0 0 0 0 0 56 104 0 3
814 752
218 752
218 749
0 1 8 0 0 0 0 0 57 105 0 4
929 761
929 993
285 993
285 747
0 1 5 0 0 0 0 0 58 87 0 4
1055 761
1055 969
337 969
337 746
0 1 25 0 0 8320 0 0 59 92 0 4
1170 761
1170 956
411 956
411 745
0 1 33 0 0 0 0 0 60 96 0 4
1277 761
1277 944
475 944
475 745
0 1 31 0 0 0 0 0 55 100 0 4
1370 761
1370 925
532 925
532 738
5 3 43 0 0 4224 0 64 65 0 0 2
1073 779
1011 779
6 1 5 0 0 0 0 64 65 0 0 2
1079 761
1011 761
5 3 44 0 0 4224 0 65 66 0 0 2
957 779
883 779
0 2 45 0 0 4096 0 0 65 108 0 5
1018 885
1018 813
1027 813
1027 770
1018 770
0 4 46 0 0 4096 0 0 65 109 0 2
987 847
987 809
5 3 47 0 0 4224 0 63 64 0 0 2
1184 779
1127 779
6 1 25 0 0 0 0 63 64 0 0 2
1190 761
1127 761
0 2 45 0 0 0 0 0 64 108 0 5
1134 885
1134 813
1143 813
1143 770
1134 770
0 4 46 0 0 0 0 0 64 109 0 2
1103 847
1103 809
5 3 48 0 0 4224 0 62 63 0 0 2
1288 779
1238 779
6 1 33 0 0 0 0 62 63 0 0 2
1294 761
1238 761
0 2 45 0 0 0 0 0 63 108 0 5
1245 885
1245 813
1254 813
1254 770
1245 770
0 4 46 0 0 0 0 0 63 109 0 2
1214 847
1214 809
6 3 49 0 0 8320 0 61 62 0 0 5
1390 756
1390 772
1363 772
1363 779
1342 779
1 5 31 0 0 0 0 62 61 0 0 6
1342 761
1376 761
1376 780
1376 780
1376 774
1384 774
0 2 45 0 0 0 0 0 62 108 0 5
1349 885
1349 813
1358 813
1358 770
1349 770
0 4 46 0 0 0 0 0 62 109 0 2
1318 847
1318 809
5 1 50 0 0 12416 0 66 61 0 0 6
829 779
826 779
826 670
1468 670
1468 756
1438 756
3 6 11 0 0 0 0 61 66 0 0 6
1438 774
1449 774
1449 712
814 712
814 761
835 761
1 6 8 0 0 0 0 66 65 0 0 2
883 761
963 761
0 2 45 0 0 0 0 0 66 108 0 5
890 885
890 813
899 813
899 770
890 770
0 4 46 0 0 0 0 0 66 109 0 2
859 847
859 809
2 1 45 0 0 20608 0 61 5 0 0 6
1445 765
1466 765
1466 825
1467 825
1467 885
705 885
1 4 46 0 0 4224 0 6 61 0 0 5
706 847
1323 847
1323 846
1414 846
1414 804
34
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
512 659 549 683
522 667 538 683
2 T1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
457 659 494 683
467 667 483 683
2 T2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
396 661 433 685
406 669 422 685
2 T3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
317 660 354 684
327 668 343 684
2 T4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
263 661 300 685
273 669 289 685
2 T5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
196 659 233 683
206 667 222 683
2 T6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
322 618 407 642
332 626 396 642
8 T States
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
415 1239 460 1263
425 1247 449 1263
3 LDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
415 1355 460 1379
425 1363 449 1379
3 ADD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
414 1484 459 1508
424 1492 448 1508
3 SUB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
413 1606 458 1630
423 1614 447 1630
3 OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
412 1731 457 1755
422 1739 446 1755
3 HLT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
606 1020 651 1044
616 1028 640 1044
3 LDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
552 1020 597 1044
562 1028 586 1044
3 ADD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
493 1019 538 1043
503 1027 527 1043
3 SUB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
432 1018 477 1042
442 1026 466 1042
3 OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
365 1015 410 1039
375 1023 399 1039
3 HLT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
451 998 552 1022
461 1006 541 1022
10 Operations
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
68 390 105 414
78 398 94 414
2 Cp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
113 389 150 413
123 397 139 413
2 Ep
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
160 388 205 412
170 396 194 412
3 Lm`
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
215 389 260 413
225 397 249 413
3 Ce`
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
344 391 389 415
354 399 378 415
3 Li`
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
398 391 443 415
408 399 432 415
3 Ei`
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
451 390 496 414
461 398 485 414
3 La`
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
507 390 544 414
517 398 533 414
2 Ea
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
669 385 706 409
679 393 695 409
2 Su
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
726 384 763 408
736 392 752 408
2 Eu
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
770 386 815 410
780 394 804 410
3 Lb`
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
820 384 865 408
830 392 854 408
3 Lo`
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
768 1324 877 1348
778 1332 866 1348
11 LDA+ADD+SUB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1026 1389 1071 1413
1036 1397 1060 1413
3 Lm`
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
985 1505 1030 1529
995 1513 1019 1529
3 Ce`
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
876 1645 921 1669
886 1653 910 1669
3 Ei`
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
