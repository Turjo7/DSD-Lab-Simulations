CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
64
13 Logic Switch~
5 37 28 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5398 0 0
2
43492.9 0
0
13 Logic Switch~
5 117 32 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7935 0 0
2
43492.9 0
0
13 Logic Switch~
5 200 32 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
356 0 0
2
43492.9 0
0
13 Logic Switch~
5 282 36 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4629 0 0
2
43492.9 0
0
13 Logic Switch~
5 126 2827 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
538 0 0
2
43492.9 0
0
13 Logic Switch~
5 232 2828 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5713 0 0
2
43492.9 0
0
13 Logic Switch~
5 342 2826 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6618 0 0
2
43492.9 0
0
2 +V
167 1193 2167 0 1 3
0 3
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3714 0 0
2
43492.9 0
0
7 Ground~
168 1071 2208 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9116 0 0
2
43492.9 0
0
5 4049~
219 37 129 0 2 22
0 4 8
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U23A
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 23 0
1 U
7960 0 0
2
43492.9 0
0
5 4049~
219 116 107 0 2 22
0 5 9
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U22F
17 -8 45 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 22 0
1 U
3886 0 0
2
43492.9 0
0
5 4049~
219 300 61 0 2 22
0 6 10
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U22E
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 22 0
1 U
3299 0 0
2
43492.9 0
0
5 4049~
219 560 26 0 2 22
0 7 11
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U22D
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 22 0
1 U
9107 0 0
2
43492.9 0
0
5 4049~
219 151 2743 0 2 22
0 14 17
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U22C
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 22 0
1 U
6556 0 0
2
43492.9 0
0
5 4049~
219 241 2737 0 2 22
0 13 16
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U22B
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 22 0
1 U
3205 0 0
2
43492.9 0
0
5 4049~
219 352 2733 0 2 22
0 12 15
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U22A
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 22 0
1 U
7255 0 0
2
43492.9 0
0
14 Logic Display~
6 1105 63 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8613 0 0
2
43492.9 0
0
14 Logic Display~
6 1058 62 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7832 0 0
2
43492.9 0
0
14 Logic Display~
6 1020 62 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8937 0 0
2
43492.9 0
0
14 Logic Display~
6 979 62 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
556 0 0
2
43492.9 0
0
5 4082~
219 486 1993 0 5 22
0 4 17 16 15 31
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U21B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 21 0
1 U
6981 0 0
2
43492.9 10
0
5 4082~
219 488 2074 0 5 22
0 8 17 16 12 30
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U21A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 21 0
1 U
8701 0 0
2
43492.9 9
0
5 4082~
219 488 2154 0 5 22
0 2 17 13 15 29
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U20B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 20 0
1 U
5540 0 0
2
43492.9 8
0
5 4082~
219 487 2231 0 5 22
0 5 17 13 12 28
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U20A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 20 0
1 U
8365 0 0
2
43492.9 7
0
5 4082~
219 488 2308 0 5 22
0 7 14 16 15 27
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U19B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 19 0
1 U
5209 0 0
2
43492.9 6
0
5 4082~
219 488 2384 0 5 22
0 5 14 16 12 26
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U19A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 19 0
1 U
3297 0 0
2
43492.9 5
0
5 4082~
219 488 2455 0 5 22
0 2 14 13 15 25
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U18B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 18 0
1 U
9904 0 0
2
43492.9 4
0
5 4082~
219 487 2537 0 5 22
0 3 14 13 12 24
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U18A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 18 0
1 U
6918 0 0
2
43492.9 3
0
8 4-In OR~
219 661 2107 0 5 22
0 31 30 29 28 23
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U17B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 17 0
1 U
7751 0 0
2
43492.9 2
0
8 4-In OR~
219 663 2415 0 5 22
0 27 26 25 24 22
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U17A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 17 0
1 U
9907 0 0
2
43492.9 1
0
5 4071~
219 831 2244 0 3 22
0 23 22 18
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 6 0
1 U
6628 0 0
2
43492.9 0
0
5 4082~
219 487 1359 0 5 22
0 5 17 16 15 41
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U16B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 16 0
1 U
4914 0 0
2
43492.9 10
0
5 4082~
219 489 1440 0 5 22
0 9 17 16 12 40
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U16A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 16 0
1 U
635 0 0
2
43492.9 9
0
5 4082~
219 489 1520 0 5 22
0 4 17 13 15 39
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U15B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 15 0
1 U
3606 0 0
2
43492.9 8
0
5 4082~
219 488 1597 0 5 22
0 6 17 13 12 38
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U15A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 15 0
1 U
8769 0 0
2
43492.9 7
0
5 4082~
219 489 1674 0 5 22
0 4 14 16 15 37
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U14B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 14 0
1 U
3887 0 0
2
43492.9 6
0
5 4082~
219 489 1750 0 5 22
0 6 14 16 12 36
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U14A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 14 0
1 U
4266 0 0
2
43492.9 5
0
5 4082~
219 489 1821 0 5 22
0 2 14 13 15 35
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U13B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 13 0
1 U
3389 0 0
2
43492.9 4
0
5 4082~
219 488 1903 0 5 22
0 3 14 13 12 34
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U13A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 13 0
1 U
8108 0 0
2
43492.9 3
0
8 4-In OR~
219 662 1473 0 5 22
0 41 40 39 38 33
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U12B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 12 0
1 U
3301 0 0
2
43492.9 2
0
8 4-In OR~
219 664 1781 0 5 22
0 37 36 35 34 32
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U12A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 12 0
1 U
3739 0 0
2
43492.9 1
0
5 4071~
219 832 1610 0 3 22
0 33 32 19
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 6 0
1 U
4610 0 0
2
43492.9 0
0
5 4082~
219 490 712 0 5 22
0 6 17 16 15 51
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U11B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 11 0
1 U
7104 0 0
2
43492.9 10
0
5 4082~
219 492 793 0 5 22
0 10 17 16 12 50
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U11A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 11 0
1 U
5233 0 0
2
43492.9 9
0
5 4082~
219 492 873 0 5 22
0 5 17 13 15 49
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U10B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
345 0 0
2
43492.9 8
0
5 4082~
219 491 950 0 5 22
0 7 17 13 12 48
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U10A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
4311 0 0
2
43492.9 7
0
5 4082~
219 492 1027 0 5 22
0 5 14 16 15 47
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U9B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 9 0
1 U
3959 0 0
2
43492.9 6
0
5 4082~
219 492 1103 0 5 22
0 7 14 16 12 46
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U9A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 9 0
1 U
9550 0 0
2
43492.9 5
0
5 4082~
219 492 1174 0 5 22
0 2 14 13 15 45
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 8 0
1 U
4183 0 0
2
43492.9 4
0
5 4082~
219 491 1256 0 5 22
0 3 14 13 12 44
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 8 0
1 U
7662 0 0
2
43492.9 3
0
8 4-In OR~
219 665 826 0 5 22
0 51 50 49 48 43
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U7B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 7 0
1 U
6373 0 0
2
43492.9 2
0
8 4-In OR~
219 667 1134 0 5 22
0 47 46 45 44 42
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
76 0 0
2
43492.9 1
0
5 4071~
219 835 963 0 3 22
0 43 42 20
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
4168 0 0
2
43492.9 0
0
5 4071~
219 835 340 0 3 22
0 53 52 21
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
9490 0 0
2
43492.9 0
0
8 4-In OR~
219 667 511 0 5 22
0 57 56 55 54 52
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U5B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
3202 0 0
2
43492.9 0
0
8 4-In OR~
219 665 203 0 5 22
0 61 60 59 58 53
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
5212 0 0
2
43492.9 0
0
5 4082~
219 491 633 0 5 22
0 3 14 13 12 54
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
5341 0 0
2
43492.9 0
0
5 4082~
219 492 551 0 5 22
0 2 14 13 15 55
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
3516 0 0
2
43492.9 0
0
5 4082~
219 492 480 0 5 22
0 4 14 16 12 56
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
6823 0 0
2
43492.9 0
0
5 4082~
219 492 404 0 5 22
0 6 14 16 15 57
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
3532 0 0
2
43492.9 0
0
5 4082~
219 491 327 0 5 22
0 2 17 13 12 58
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
3978 0 0
2
43492.9 0
0
5 4082~
219 492 250 0 5 22
0 6 17 13 15 59
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
4691 0 0
2
43492.9 0
0
5 4082~
219 492 170 0 5 22
0 11 17 16 12 60
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 1 0
1 U
5392 0 0
2
43492.9 0
0
5 4082~
219 490 89 0 5 22
0 7 17 16 15 61
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
3264 0 0
2
43492.9 0
0
179
0 1 3 0 0 8192 0 0 28 4 0 5
1175 2176
1175 2504
385 2504
385 2524
463 2524
0 1 3 0 0 0 0 0 39 4 0 6
1152 2081
1122 2081
1122 1869
439 1869
439 1890
464 1890
0 1 3 0 0 8192 0 0 50 4 0 6
1152 2142
1108 2142
1108 1206
406 1206
406 1243
467 1243
1 1 3 0 0 8320 0 8 57 0 0 6
1193 2176
1152 2176
1152 596
426 596
426 620
467 620
0 1 2 0 0 12288 0 0 27 21 0 6
1071 2190
995 2190
995 2490
423 2490
423 2442
464 2442
0 1 2 0 0 0 0 0 38 21 0 5
997 2180
997 1855
439 1855
439 1808
465 1808
0 1 2 0 0 4096 0 0 49 21 0 7
1034 2180
1034 1194
536 1194
536 1140
451 1140
451 1161
468 1161
0 1 2 0 0 4096 0 0 58 21 0 5
1011 2180
1011 583
446 583
446 538
468 538
0 1 4 0 0 4096 0 0 59 14 0 6
14 196
565 196
565 438
438 438
438 467
468 467
0 1 5 0 0 4224 0 0 26 34 0 3
137 32
137 2371
464 2371
0 1 6 0 0 8320 0 0 37 35 0 4
232 49
199 49
199 1737
465 1737
0 1 7 0 0 4096 0 0 48 36 0 3
349 36
349 1090
468 1090
0 1 7 0 0 12416 0 0 25 32 0 7
495 26
495 5
899 5
899 2267
446 2267
446 2295
464 2295
0 1 4 0 0 8192 0 0 36 33 0 4
71 54
14 54
14 1661
465 1661
0 1 5 0 0 0 0 0 47 34 0 3
162 32
162 1014
468 1014
0 1 6 0 0 0 0 0 60 35 0 4
232 97
217 97
217 391
468 391
0 1 2 0 0 4224 0 0 61 21 0 5
1051 2180
1051 281
444 281
444 314
467 314
0 1 5 0 0 128 0 0 24 34 0 3
148 32
148 2218
463 2218
0 1 6 0 0 128 0 0 35 35 0 4
232 39
255 39
255 1584
464 1584
0 1 7 0 0 128 0 0 46 36 0 3
405 36
405 937
467 937
1 1 2 0 0 128 0 9 23 0 0 5
1071 2202
1071 2180
413 2180
413 2141
464 2141
0 1 4 0 0 0 0 0 34 33 0 4
71 40
88 40
88 1507
465 1507
0 1 5 0 0 0 0 0 45 34 0 4
173 45
193 45
193 860
468 860
0 1 6 0 0 0 0 0 62 30 0 3
270 61
270 237
468 237
2 1 8 0 0 4224 0 10 22 0 0 3
40 147
40 2061
464 2061
2 1 9 0 0 4224 0 11 33 0 0 3
119 125
119 1427
465 1427
0 1 4 0 0 0 0 0 10 33 0 3
71 66
40 66
40 111
0 1 5 0 0 0 0 0 11 34 0 3
173 54
119 54
119 89
2 1 10 0 0 8320 0 12 44 0 0 4
321 61
337 61
337 780
468 780
0 1 6 0 0 0 0 0 12 35 0 3
232 63
232 61
285 61
2 1 11 0 0 12416 0 13 63 0 0 6
581 26
602 26
602 130
444 130
444 157
468 157
0 1 7 0 0 128 0 0 13 36 0 3
379 36
379 26
545 26
1 1 4 0 0 8320 0 1 21 0 0 4
49 28
71 28
71 1980
462 1980
1 1 5 0 0 128 0 2 32 0 0 4
129 32
173 32
173 1346
463 1346
1 1 6 0 0 128 0 3 43 0 0 4
212 32
232 32
232 699
466 699
1 1 7 0 0 128 0 4 64 0 0 4
294 36
460 36
460 76
466 76
0 4 12 0 0 8192 0 0 28 112 0 3
310 2552
310 2551
463 2551
0 4 12 0 0 8192 0 0 39 112 0 3
310 1915
310 1917
464 1917
0 4 12 0 0 4096 0 0 50 112 0 2
310 1270
467 1270
0 4 12 0 0 0 0 0 57 112 0 3
310 648
310 647
467 647
0 3 13 0 0 8192 0 0 28 104 0 3
206 2541
206 2542
463 2542
0 3 13 0 0 4096 0 0 39 104 0 2
206 1908
464 1908
0 3 13 0 0 4096 0 0 50 104 0 2
206 1261
467 1261
0 3 13 0 0 0 0 0 57 104 0 2
206 638
467 638
0 2 14 0 0 8192 0 0 28 84 0 3
103 2530
103 2533
463 2533
0 2 14 0 0 8192 0 0 39 84 0 3
103 1901
103 1899
464 1899
0 2 14 0 0 8192 0 0 50 84 0 3
103 1253
103 1252
467 1252
0 2 14 0 0 0 0 0 57 84 0 3
103 630
103 629
467 629
0 4 15 0 0 8192 0 0 27 127 0 3
355 2468
355 2469
464 2469
0 4 15 0 0 4096 0 0 38 127 0 2
355 1835
465 1835
0 4 15 0 0 8192 0 0 49 127 0 3
355 1190
355 1188
468 1188
0 4 15 0 0 0 0 0 58 127 0 3
355 566
355 565
468 565
0 3 13 0 0 0 0 0 27 104 0 3
206 2459
206 2460
464 2460
0 3 13 0 0 0 0 0 38 104 0 3
206 1827
206 1826
465 1826
0 3 13 0 0 8192 0 0 49 104 0 3
206 1177
206 1179
468 1179
0 3 13 0 0 0 0 0 58 104 0 3
206 554
206 556
468 556
0 2 14 0 0 0 0 0 27 84 0 3
103 2453
103 2451
464 2451
0 2 14 0 0 0 0 0 38 84 0 3
103 1816
103 1817
465 1817
0 2 14 0 0 8192 0 0 49 84 0 3
103 1172
103 1170
468 1170
0 2 14 0 0 0 0 0 58 84 0 3
103 546
103 547
468 547
0 4 12 0 0 0 0 0 26 112 0 3
310 2400
310 2398
464 2398
0 4 12 0 0 0 0 0 37 112 0 3
310 1765
310 1764
465 1764
0 4 12 0 0 8192 0 0 48 112 0 3
310 1118
310 1117
468 1117
0 4 12 0 0 0 0 0 59 112 0 3
310 495
310 494
468 494
0 3 16 0 0 8192 0 0 26 128 0 3
244 2388
244 2389
464 2389
0 3 16 0 0 8192 0 0 37 128 0 3
244 1757
244 1755
465 1755
0 3 16 0 0 4096 0 0 48 128 0 2
244 1108
468 1108
0 3 16 0 0 0 0 0 59 128 0 3
244 484
244 485
468 485
0 2 14 0 0 0 0 0 26 84 0 2
103 2380
464 2380
0 2 14 0 0 0 0 0 37 84 0 3
103 1748
103 1746
465 1746
0 2 14 0 0 0 0 0 48 84 0 3
103 1101
103 1099
468 1099
0 2 14 0 0 0 0 0 59 84 0 3
103 474
103 476
468 476
0 4 15 0 0 0 0 0 25 127 0 3
355 2323
355 2322
464 2322
0 4 15 0 0 0 0 0 36 127 0 2
355 1688
465 1688
0 4 15 0 0 0 0 0 47 127 0 2
355 1041
468 1041
0 4 15 0 0 0 0 0 60 127 0 3
355 417
355 418
468 418
0 3 16 0 0 0 0 0 25 128 0 3
244 2314
244 2313
464 2313
0 3 16 0 0 0 0 0 36 128 0 3
244 1680
244 1679
465 1679
0 3 16 0 0 0 0 0 47 128 0 3
244 1033
244 1032
468 1032
0 3 16 0 0 0 0 0 60 128 0 3
244 408
244 409
468 409
0 2 14 0 0 0 0 0 25 84 0 3
103 2303
103 2304
464 2304
0 2 14 0 0 0 0 0 36 84 0 2
103 1670
465 1670
0 2 14 0 0 0 0 0 47 84 0 3
103 1024
103 1023
468 1023
0 2 14 0 0 8320 0 0 60 133 0 4
166 2780
103 2780
103 400
468 400
0 4 12 0 0 0 0 0 24 112 0 2
310 2245
463 2245
0 4 12 0 0 0 0 0 35 112 0 2
310 1611
464 1611
0 4 12 0 0 0 0 0 46 112 0 2
310 964
467 964
0 4 12 0 0 0 0 0 61 112 0 2
310 341
467 341
0 3 13 0 0 0 0 0 24 104 0 3
206 2235
206 2236
463 2236
0 3 13 0 0 0 0 0 35 104 0 3
206 1600
206 1602
464 1602
0 3 13 0 0 0 0 0 46 104 0 2
206 955
467 955
0 3 13 0 0 0 0 0 61 104 0 3
206 331
206 332
467 332
0 2 17 0 0 8192 0 0 24 132 0 3
154 2225
154 2227
463 2227
0 2 17 0 0 8192 0 0 35 132 0 3
154 1590
154 1593
464 1593
0 2 17 0 0 8192 0 0 46 132 0 3
154 947
154 946
467 946
0 2 17 0 0 0 0 0 61 132 0 3
154 324
154 323
467 323
0 4 15 0 0 0 0 0 23 127 0 3
355 2167
355 2168
464 2168
0 4 15 0 0 0 0 0 34 127 0 3
355 1533
355 1534
465 1534
0 4 15 0 0 0 0 0 45 127 0 3
355 888
355 887
468 887
0 4 15 0 0 0 0 0 62 127 0 3
355 263
355 264
468 264
0 3 13 0 0 0 0 0 23 104 0 3
206 2156
206 2159
464 2159
0 3 13 0 0 0 0 0 34 104 0 2
206 1525
465 1525
0 3 13 0 0 0 0 0 45 104 0 2
206 878
468 878
0 3 13 0 0 8320 0 0 62 134 0 4
264 2774
206 2774
206 255
468 255
0 2 17 0 0 0 0 0 23 132 0 3
154 2148
154 2150
464 2150
0 2 17 0 0 0 0 0 34 132 0 3
154 1515
154 1516
465 1516
0 2 17 0 0 8192 0 0 45 132 0 3
154 868
154 869
468 869
0 2 17 0 0 0 0 0 62 132 0 3
154 245
154 246
468 246
0 4 12 0 0 0 0 0 22 112 0 2
310 2088
464 2088
0 4 12 0 0 0 0 0 33 112 0 3
310 1455
310 1454
465 1454
0 4 12 0 0 0 0 0 44 112 0 3
310 805
310 807
468 807
0 4 12 0 0 8320 0 0 63 135 0 4
365 2770
310 2770
310 184
468 184
0 3 16 0 0 0 0 0 22 128 0 3
244 2078
244 2079
464 2079
0 2 17 0 0 0 0 0 22 132 0 3
154 2071
154 2070
464 2070
0 3 16 0 0 0 0 0 33 128 0 3
244 1443
244 1445
465 1445
0 2 17 0 0 0 0 0 33 132 0 2
154 1436
465 1436
0 3 16 0 0 0 0 0 44 128 0 3
244 800
244 798
468 798
0 2 17 0 0 0 0 0 44 132 0 3
154 787
154 789
468 789
0 3 16 0 0 0 0 0 63 128 0 3
244 174
244 175
468 175
0 2 17 0 0 0 0 0 63 132 0 3
154 165
154 166
468 166
0 4 15 0 0 0 0 0 21 127 0 3
355 2008
355 2007
462 2007
0 3 16 0 0 0 0 0 21 128 0 3
244 1999
244 1998
462 1998
0 4 15 0 0 0 0 0 32 127 0 3
355 1374
355 1373
463 1373
0 3 16 0 0 0 0 0 32 128 0 3
244 1365
244 1364
463 1364
0 4 15 0 0 0 0 0 43 127 0 3
355 724
355 726
466 726
0 3 16 0 0 0 0 0 43 128 0 3
244 715
244 717
466 717
2 4 15 0 0 4224 0 16 64 0 0 3
355 2715
355 103
466 103
2 3 16 0 0 4224 0 15 64 0 0 3
244 2719
244 94
466 94
0 2 17 0 0 0 0 0 21 132 0 3
154 1987
154 1989
462 1989
0 2 17 0 0 0 0 0 32 132 0 4
154 1350
438 1350
438 1355
463 1355
0 2 17 0 0 0 0 0 43 132 0 3
154 706
154 708
466 708
2 2 17 0 0 4224 0 14 64 0 0 3
154 2725
154 85
466 85
1 1 14 0 0 0 0 5 14 0 0 5
138 2827
166 2827
166 2767
154 2767
154 2761
1 1 13 0 0 0 0 6 15 0 0 5
244 2828
264 2828
264 2766
244 2766
244 2755
1 1 12 0 0 0 0 7 16 0 0 5
354 2826
365 2826
365 2765
355 2765
355 2751
3 1 18 0 0 8320 0 31 20 0 0 3
864 2244
979 2244
979 80
3 1 19 0 0 8320 0 42 19 0 0 5
865 1610
968 1610
968 107
1020 107
1020 80
3 1 20 0 0 8320 0 53 18 0 0 5
868 963
1034 963
1034 121
1058 121
1058 80
3 1 21 0 0 8320 0 54 17 0 0 3
868 340
1105 340
1105 81
5 2 22 0 0 8336 0 30 31 0 0 4
696 2415
774 2415
774 2253
818 2253
5 1 23 0 0 8336 0 29 31 0 0 4
694 2107
773 2107
773 2235
818 2235
5 4 24 0 0 4240 0 28 30 0 0 4
508 2537
628 2537
628 2429
646 2429
5 3 25 0 0 4240 0 27 30 0 0 4
509 2455
618 2455
618 2420
646 2420
5 2 26 0 0 4240 0 26 30 0 0 4
509 2384
617 2384
617 2411
646 2411
5 1 27 0 0 4240 0 25 30 0 0 4
509 2308
629 2308
629 2402
646 2402
5 4 28 0 0 4240 0 24 29 0 0 4
508 2231
630 2231
630 2121
644 2121
5 3 29 0 0 4240 0 23 29 0 0 4
509 2154
603 2154
603 2112
644 2112
5 2 30 0 0 4240 0 22 29 0 0 4
509 2074
603 2074
603 2103
644 2103
5 1 31 0 0 4240 0 21 29 0 0 4
507 1993
629 1993
629 2094
644 2094
5 2 32 0 0 8320 0 41 42 0 0 4
697 1781
775 1781
775 1619
819 1619
5 1 33 0 0 8320 0 40 42 0 0 4
695 1473
774 1473
774 1601
819 1601
5 4 34 0 0 4224 0 39 41 0 0 4
509 1903
629 1903
629 1795
647 1795
5 3 35 0 0 4224 0 38 41 0 0 4
510 1821
619 1821
619 1786
647 1786
5 2 36 0 0 4224 0 37 41 0 0 4
510 1750
618 1750
618 1777
647 1777
5 1 37 0 0 4224 0 36 41 0 0 4
510 1674
630 1674
630 1768
647 1768
5 4 38 0 0 4224 0 35 40 0 0 4
509 1597
631 1597
631 1487
645 1487
5 3 39 0 0 4224 0 34 40 0 0 4
510 1520
604 1520
604 1478
645 1478
5 2 40 0 0 4224 0 33 40 0 0 4
510 1440
604 1440
604 1469
645 1469
5 1 41 0 0 4224 0 32 40 0 0 4
508 1359
630 1359
630 1460
645 1460
5 2 42 0 0 8320 0 52 53 0 0 4
700 1134
778 1134
778 972
822 972
5 1 43 0 0 8320 0 51 53 0 0 4
698 826
777 826
777 954
822 954
5 4 44 0 0 4224 0 50 52 0 0 4
512 1256
632 1256
632 1148
650 1148
5 3 45 0 0 4224 0 49 52 0 0 4
513 1174
622 1174
622 1139
650 1139
5 2 46 0 0 4224 0 48 52 0 0 4
513 1103
621 1103
621 1130
650 1130
5 1 47 0 0 4224 0 47 52 0 0 4
513 1027
633 1027
633 1121
650 1121
5 4 48 0 0 4224 0 46 51 0 0 4
512 950
634 950
634 840
648 840
5 3 49 0 0 4224 0 45 51 0 0 4
513 873
607 873
607 831
648 831
5 2 50 0 0 4224 0 44 51 0 0 4
513 793
607 793
607 822
648 822
5 1 51 0 0 4224 0 43 51 0 0 4
511 712
633 712
633 813
648 813
5 2 52 0 0 8320 0 55 54 0 0 4
700 511
778 511
778 349
822 349
5 1 53 0 0 8320 0 56 54 0 0 4
698 203
777 203
777 331
822 331
5 4 54 0 0 4224 0 57 55 0 0 4
512 633
632 633
632 525
650 525
5 3 55 0 0 4224 0 58 55 0 0 4
513 551
622 551
622 516
650 516
5 2 56 0 0 4224 0 59 55 0 0 4
513 480
621 480
621 507
650 507
5 1 57 0 0 4224 0 60 55 0 0 4
513 404
633 404
633 498
650 498
5 4 58 0 0 4224 0 61 56 0 0 4
512 327
634 327
634 217
648 217
5 3 59 0 0 4224 0 62 56 0 0 4
513 250
607 250
607 208
648 208
5 2 60 0 0 4224 0 63 56 0 0 4
513 170
607 170
607 199
648 199
5 1 61 0 0 4224 0 64 56 0 0 4
511 89
633 89
633 190
648 190
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
