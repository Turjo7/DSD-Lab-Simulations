CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 40 30 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9961490 0
0
6 Title:
5 Name:
0
0
0
16
5 4071~
219 901 608 0 1 22
0 0
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
5130 0 0
2
43513.9 0
0
5 4049~
219 608 618 0 1 22
0 0
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
391 0 0
2
43513.9 0
0
5 4073~
219 813 594 0 1 22
0 0
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
3124 0 0
2
43513.9 0
0
5 4030~
219 682 545 0 1 22
0 0
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
3421 0 0
2
43513.9 0
0
13 Logic Switch~
5 696 404 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8157 0 0
2
43513.9 0
0
13 Logic Switch~
5 413 414 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 S2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5572 0 0
2
43513.9 0
0
13 Logic Switch~
5 513 417 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8901 0 0
2
43513.9 0
0
13 Logic Switch~
5 592 418 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7361 0 0
2
43513.9 0
0
13 Logic Switch~
5 141 199 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4747 0 0
2
43513.9 0
0
13 Logic Switch~
5 256 200 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
972 0 0
2
43513.9 0
0
13 Logic Switch~
5 365 202 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3472 0 0
2
43513.9 0
0
13 Logic Switch~
5 476 200 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9998 0 0
2
43513.9 0
0
13 Logic Switch~
5 136 90 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3536 0 0
2
43513.9 0
0
13 Logic Switch~
5 254 94 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4597 0 0
2
43513.9 0
0
13 Logic Switch~
5 370 94 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3835 0 0
2
43513.9 0
0
13 Logic Switch~
5 472 92 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3670 0 0
2
43513.9 0
0
8
1 2 0 0 0 0 0 16 1 0 0 4
484 92
842 92
842 617
888 617
4 1 0 0 0 0 0 3 1 0 0 4
834 594
862 594
862 599
888 599
2 3 0 0 0 0 0 2 3 0 0 4
629 618
761 618
761 603
789 603
1 1 0 0 0 0 0 8 2 0 0 6
604 418
618 418
618 577
571 577
571 618
593 618
1 2 0 0 0 0 0 6 3 0 0 4
425 414
451 414
451 594
789 594
3 1 0 0 0 0 0 4 3 0 0 4
715 545
760 545
760 585
789 585
1 2 0 0 0 0 0 12 4 0 0 6
488 200
515 200
515 355
375 355
375 554
666 554
1 1 0 0 0 0 0 7 4 0 0 4
525 417
547 417
547 536
666 536
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
889 592 926 616
899 600 915 616
2 X0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
